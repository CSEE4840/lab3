0F
30
40
47
88
90
90
90
FF
00
00
FF
00
00
00
00
FF
00
00
E0
10
08
08
08
FF
00
00
07
08
10
10
10
F0
0C
02
E2
11
09
09
09
09
09
09
11
E2
02
0C
F0
00
00
00
00
FF
00
00
00
00
00
00
07
08
10
10
10
00
00
00
E0
10
08
08
08
90
90
90
90
90
90
90
90
00
00
00
18
18
00
00
00
08
08
08
08
08
08
08
08
10
10
10
10
10
10
10
10
09
09
09
09
09
09
09
09
09
09
09
11
E1
01
01
01
90
90
90
88
87
80
80
80
00
00
00
FF
00
00
00
00
10
10
10
08
07
00
00
00
08
08
08
10
E0
00
00
00
90
90
90
88
47
40
30
0F
3C
7E
FF
FF
FF
FF
7E
3C
08
08
08
04
03
00
00
00
10
10
10
20
C0
00
00
00
00
00
00
00
0F
08
08
09
00
00
00
00
FF
01
01
FF
00
00
00
00
FF
80
80
FF
00
00
00
00
F0
10
10
90
00
00
00
00
03
04
08
08
00
00
00
00
FF
00
00
FF
00
00
00
00
C0
20
10
10
09
08
08
0F
00
00
00
00
00
00
00
00
00
FF
FF
00
90
10
10
F0
00
00
00
00
08
08
04
03
00
00
00
00
10
10
20
C0
00
00
00
00
80
80
80
87
88
90
90
90
01
01
01
E1
11
09
09
09
00
00
00
00
00
00
00
00