// left
0000
0000
07c0
1ff0
3ff8
3ff8
0ffc
03fc
00fc
03fc
0ffc
3ff8
3ff8
1ff0
07c0
0000




// up
0000
0000
0c30
1c1c
1e3c
3e3e
3f7e
3ffe
3ffe
1ffc
1ffc
0ff8
03e0
0000
0000


// down
0000
0000
0000
03e0
0ff8
1ffc
1ffc
3ffe
3ffe
3f7e
3e3e
1e3c
1c1c
0c30
0000
0000



// right
0000
0000
03e0
0ff8
1ffc
1ffc
3ff0
3fc0
3f00
3fc0
3ff0
1ffc
1ffc
0ff8
03e0
0000



//eat
0000
0000
03e0
0ff8
1ffc
1ffc
3ffe
3ffe
3ffe
3ffe
3ffe
1ffc
1ffc
0ff8
03e0
0000


07E0  
0000  
0000  

