0000
07C0
1FF0
3FF8
3FF8
0FFC
01FC
00FC
01FC
1FFC
3FF8
3FF8
1FF0
07C0
0000
0000
