// left
assign pacman_left[0] = 16'h0000;
assign pacman_left[1] = 16'h07C0;
assign pacman_left[2] = 16'h1FF0;
assign pacman_left[3] = 16'h3FF8;
assign pacman_left[4] = 16'h3FF8;
assign pacman_left[5] = 16'h0FFC;
assign pacman_left[6] = 16'h01FC;
assign pacman_left[7] = 16'h00FC;
assign pacman_left[8] = 16'h01FC;
assign pacman_left[9] = 16'h1FFC;
assign pacman_left[10] = 16'h3FF8;
assign pacman_left[11] = 16'h3FF8;
assign pacman_left[12] = 16'h1FF0;
assign pacman_left[13] = 16'h07C0;
assign pacman_left[14] = 16'h0000;
assign pacman_left[15] = 16'h0000;

// up
assign pacman_up[0] = 16'h0000;
assign pacman_up[1] = 16'h0000;
assign pacman_up[2] = 16'h1830;
assign pacman_up[3] = 16'h3878;
assign pacman_up[4] = 16'h3C78;
assign pacman_up[5] = 16'h7C7C;
assign pacman_up[6] = 16'h7C7C;
assign pacman_up[7] = 16'h7EFC;
assign pacman_up[8] = 16'h7FFC;
assign pacman_up[9] = 16'h7FFC;
assign pacman_up[10] = 16'h3FF8;
assign pacman_up[11] = 16'h3FF0;
assign pacman_up[12] = 16'h1FC0;
assign pacman_up[13] = 16'h07C0;
assign pacman_up[14] = 16'h0000;
assign pacman_up[15] = 16'h0000;

// down
assign pacman_down[0] = 16'h0000;
assign pacman_down[1] = 16'h0000;
assign pacman_down[2] = 16'h07C0;
assign pacman_down[3] = 16'h1FE0;
assign pacman_down[4] = 16'h3FF0;
assign pacman_down[5] = 16'h3FF8;
assign pacman_down[6] = 16'h7FFC;
assign pacman_down[7] = 16'h7FFC;
assign pacman_down[8] = 16'h7EFC;
assign pacman_down[9] = 16'h7C7C;
assign pacman_down[10] = 16'h7C7C;
assign pacman_down[11] = 16'h3C78;
assign pacman_down[12] = 16'h3878;
assign pacman_down[13] = 16'h1830;
assign pacman_down[14] = 16'h0000;
assign pacman_down[15] = 16'h0000;

// right
assign pacman_right[0] = 16'h0000;
assign pacman_right[1] = 16'h03E0;
assign pacman_right[2] = 16'h0FF8;
assign pacman_right[3] = 16'h1FFC;
assign pacman_right[4] = 16'h1FFC;
assign pacman_right[5] = 16'h3F80;
assign pacman_right[6] = 16'h3F00;
assign pacman_right[7] = 16'h3F80;
assign pacman_right[8] = 16'h3FF0;
assign pacman_right[9] = 16'h3FF8;
assign pacman_right[10] = 16'h1FFC;
assign pacman_right[11] = 16'h0FFC;
assign pacman_right[12] = 16'h07F8;
assign pacman_right[13] = 16'h03E0;
assign pacman_right[14] = 16'h0000;
assign pacman_right[15] = 16'h0000;
