localparam logic [1:0] GHOST_DOWN [0:15][0:15] = '{
'{0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0},
'{0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0},
'{0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0},
'{0,0,1,1,2,2,1,1,2,2,1,1,1,0,0,0},
'{0,0,1,2,2,2,2,1,2,2,2,2,1,0,0,0},
'{0,0,1,2,2,2,2,1,2,2,2,2,1,0,0,0},
'{0,1,1,2,3,3,2,1,2,3,3,2,1,1,0,0},
'{0,1,1,1,3,3,1,1,1,3,3,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,0,1,1,1,0,0,1,1,1,0,1,1,0},
'{0,1,0,0,0,1,1,0,0,1,1,0,0,0,1,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
};
