00000000
00003C00
00FFFF00
03FFFFC0
114719DC
1CBAAE1C
1CBAAE1C
72B29CF6
74F33DFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
6E1C3B1A
43198642
00000000
