18
3C
66
C3
C3
FF
C3
C3
C3
C3
00
00
00
00
00
00
FE
66
66
66
7C
66
66
66
66
FE
00
00
00
00
00
00
3C
66
C2
C0
C0
C0
C0
C2
66
3C
00
00
00
00
00
00
FC
66
63
63
63
63
63
63
66
FC
00
00
00
00
00
00
FF
63
68
68
78
68
68
60
63
FF
00
00
00
00
00
00
FF
63
68
68
78
68
68
60
60
F0
00
00
00
00
00
00
3C
66
C2
C0
C0
CF
C3
C3
66
3C
00
00
00
00
00
00
C3
C3
C3
C3
FF
C3
C3
C3
C3
C3
00
00
00
00
00
00
3C
18
18
18
18
18
18
18
18
3C
00
00
00
00
00
00
1F
0C
0C
0C
0C
0C
CC
CC
78
30
00
00
00
00
00
00
E7
66
6C
78
70
78
6C
66
66
E7
00
00
00
00
00
00
F0
60
60
60
60
60
63
63
63
FF
00
00
00
00
00
00
C3
E7
FF
DB
C3
C3
C3
C3
C3
C3
00
00
00
00
00
00
C3
E3
F3
DB
CF
C7
C3
C3
C3
C3
00
00
00
00
00
00
3C
66
C3
C3
C3
C3
C3
C3
66
3C
00
00
00
00
00
00
FE
66
66
66
7E
60
60
60
60
F0
00
00
00
00
00
00
3C
66
C3
C3
C3
C3
CB
C7
66
3F
00
00
00
00
00
00
FE
66
66
66
7C
78
6C
66
66
E7
00
00
00
00
00
00
3E
66
C0
C0
7C
06
03
C3
66
3C
00
00
00
00
00
00
FF
DB
99
18
18
18
18
18
18
3C
00
00
00
00
00
00
C3
C3
C3
C3
C3
C3
C3
C3
66
3C
00
00
00
00
00
00
C3
C3
C3
C3
C3
C3
66
3C
18
18
00
00
00
00
00
00
C3
C3
C3
C3
C3
DB
FF
E7
C3
C3
00
00
00
00
00
00
C3
66
3C
18
18
3C
66
C3
C3
C3
00
00
00
00
00
00
C3
C3
66
3C
18
18
18
18
18
3C
00
00
00
00
00
00
FF
06
0C
18
30
60
C0
C0
C3
FF
00
00
00
00
00
00
3C
66
C3
C7
CF
DB
E3
C3
66
3C
00
00
00
00
00
00
18
38
78
18
18
18
18
18
18
7E
00
00
00
00
00
00
3C
66
C3
03
06
0C
18
30
60
FF
00
00
00
00
00
00
3C
66
C3
03
1E
03
03
C3
66
3C
00
00
00
00
00
00
06
0E
1E
36
66
FF
06
06
06
0F
00
00
00
00
00
00
FF
C0
C0
FC
06
03
03
C3
66
3C
00
00
00
00
00
00
3C
66
C0
C0
FC
C3
C3
C3
66
3C
00
00
00
00
00
00
FF
03
06
0C
18
30
60
60
60
60
00
00
00
00
00
00
3C
66
C3
66
3C
66
C3
C3
66
3C
00
00
00
00
00
00
3C
66
C3
C3
67
3F
03
03
66
3C
00
00
00
00
00
00
