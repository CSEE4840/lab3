2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h2 2'h2 2'h2 2'h2 2'h2 2'h1 2'h2 2'h2 2'h2 2'h2 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h0 2'h0 2'h0
2'h0 2'h1 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h0 2'h1 2'h1 2'h1 2'h0 2'h0 2'h1 2'h1 2'h1 2'h0 2'h1 2'h1 2'h0
2'h0 2'h1 2'h0 2'h0 2'h0 2'h1 2'h1 2'h0 2'h0 2'h1 2'h1 2'h0 2'h0 2'h0 2'h1 2'h0
2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0

0000000000000000
0000001111000000
0000111111110000
0001111111111000
0011122111221100
0011222212222100
0011223312233100
0111223312233110
0111122111221110
0111111111111110
0111111111111110
0111111111111110
0111111111111110
0110111001110110
0100011001100010
0000000000000000
