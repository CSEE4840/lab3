reg [15:0] pacman_left [0:15] = '{
    16'b0000000000000000,
    16'b0000011111000000,
    16'b0001111111110000,
    16'b0011111111111000,
    16'b0011111111111000,
    16'b0000111111111100,
    16'b0000000111111100,
    16'b0000000011111100,
    16'b0000000111111100,
    16'b0001111111111100,
    16'b0011111111111000,
    16'b0011111111111000,
    16'b0001111111110000,
    16'b0000011111000000,
    16'b0000000000000000,
    16'b0000000000000000
};

reg [15:0] pacman_up [0:15] = '{
    16'b0000000000000000,
    16'b0000000000000000,
    16'b0001100000110000,
    16'b0011100001111000,
    16'b0011110001111000,
    16'b0111110001111100,
    16'b0111110001111100,
    16'b0111111011111100,
    16'b0111111111111100,
    16'b0111111111111100,
    16'b0011111111111000,
    16'b0011111111110000,
    16'b0001111111000000,
    16'b0000011111000000,
    16'b0000000000000000,
    16'b0000000000000000
};

reg [15:0] pacman_right [0:15] = '{
    16'b0000000000000000,
    16'b0000001111100000,
    16'b0000111111111000,
    16'b0001111111111100,
    16'b0001111111111100,
    16'b0011111110000000,
    16'b0011111100000000,
    16'b0011111110000000,
    16'b0011111111110000,
    16'b0011111111111000,
    16'b0001111111111100,
    16'b0000111111111100,
    16'b0000011111111000,
    16'b0000001111100000,
    16'b0000000000000000,
    16'b0000000000000000
};

reg [15:0] pacman_down [0:15] = '{
    16'b0000000000000000,
    16'b0000000000000000,
    16'b0000011111000000,
    16'b0001111111100000,
    16'b0011111111110000,
    16'b0011111111111000,
    16'b0111111111111100,
    16'b0111111111111100,
    16'b0111111011111100,
    16'b0111110001111100,
    16'b0111110001111100,
    16'b0011110001111000,
    16'b0011100001111000,
    16'b0001100000110000,
    16'b0000000000000000,
    16'b0000000000000000
};
