00000000
00003C00
00FFFF00
03FFFFC0
114719DC
1CBAAE1C
1DCECE1C
73CECE7E
74719DFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
6E1C3B1A
43198642
00000000


localparam logic [1:0] GHOST_LEFT [0:15][0:15] = '{
'{0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0},
'{0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0},
'{0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0},
'{0,0,1,1,2,2,1,1,2,2,1,1,1,0,0,0},
'{0,0,1,2,2,2,2,1,2,2,2,2,1,0,0,0},
'{0,0,1,3,3,2,2,1,3,3,2,2,1,0,0,0},
'{0,1,1,3,3,2,2,1,3,3,2,2,1,1,0,0},
'{0,1,1,1,2,2,1,1,2,2,1,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0},
'{0,1,1,0,1,1,1,0,0,1,1,1,0,1,1,0},
'{0,1,0,0,0,1,1,0,0,1,1,0,0,0,1,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
};
