// left
0000
0000
07E0
0FFF
1FFF
1FFF
03FF
00FF
001F
00FF
03FF
1FFF
1FFF
0FFF
07E0
0000



// up
0000
0000
0C30
1C0E
1E3E
3E3F
3F7F
3FFF
3FFF
1FFE
1FFE
0FFC
03E0
0000
0000


// down
0000
0000
0000
03E0
0FFC
1FFE
1FFE
3FFF
3FFF
3F7F
3E3F
1E3E
1C0E
0C30
0000
0000


// right
0000
0000
03E0
0FFC
1FFE
1FFE
1FF0
0FF0
07E0
0FF0
1FF0
1FFE
1FFE
0FFC
03E0
0000


//eat
0000
0000
03E0
0FFC
1FFE
1FFE
3FFF
3FFF
3FFF
3FFF
3FFF
1FFE
1FFE
0FFC
03E0
0000

07E0  
0000  
0000  

