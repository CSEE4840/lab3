module vga_ball (
    input clk,
    input reset,
    input [15:0] writedata,
    input write,
    input chipselect,
    input [2:0] address,

    output reg [7:0] VGA_R, VGA_G, VGA_B,
    output VGA_CLK, VGA_HS, VGA_VS,
    output VGA_BLANK_n, VGA_SYNC_n
);

    // VGA sync counters
    wire [10:0] hcount;
    wire [9:0]  vcount;

    wire [6:0] tile_x = hcount[10:3];
    wire [5:0] tile_y = vcount[9:3];
    wire [2:0] tx = hcount[2:0];
    wire [2:0] ty = vcount[2:0];

    wire [5:0] tile_id = tiles[tile_y * 80 + tile_x];
    // VGA sync generator instance
    vga_counters counters_inst (
        .clk50(clk),
        .hcount(hcount),
        .vcount(vcount),
        .VGA_CLK(VGA_CLK),
        .VGA_HS(VGA_HS),
        .VGA_VS(VGA_VS),
        .VGA_BLANK_n(VGA_BLANK_n),
        .VGA_SYNC_n(VGA_SYNC_n)
    );

    // Tile memory (4800 tiles, each stores 6 bits for tile ID)
    reg [5:0] tiles [0:4799];

    // Tile bitmaps (41 tile types, each 8 rows of 8 bits)
    logic [7:0] tile_bitmaps [0:39][0:7] = '{
        '{8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000},
        '{8'b00000000,8'b00000000,8'b00011000,8'b00011000,8'b00011000,8'b00011000,8'b00000000,8'b00000000},
        '{8'b11111100,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000},
        '{8'b00111111,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011},
        '{8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11111100},
        '{8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00111111},
        '{8'b11111111,8'b00000000,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100},
        '{8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00000000,8'b11111111},
        '{8'b11000000,8'b11000000,8'b11000000,8'b11111111,8'b11111111,8'b11000000,8'b11000000,8'b11000000},
        '{8'b00000011,8'b00000011,8'b00000011,8'b11111111,8'b11111111,8'b00000011,8'b00000011,8'b00000011},
        '{8'b00111100,8'b00111100,8'b00111100,8'b11111111,8'b11111111,8'b00111100,8'b00111100,8'b00111100},
        '{8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111},
        '{8'b11111111,8'b11111111,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000},
        '{8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b11111111,8'b11111111},
        '{8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000},
        '{8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011},
        '{8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b11111111},
        '{8'b00000000,8'b00000000,8'b11111111,8'b11111111,8'b00000000,8'b00000000,8'b00000000,8'b00000000},
        '{8'b00110000,8'b00110000,8'b00110000,8'b00110000,8'b00110000,8'b00110000,8'b00110000,8'b00110000},
        '{8'b11111111,8'b11111111,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000},
        '{8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b11111111,8'b11111111},
        '{8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000},
        '{8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011},
        '{8'b00000000,8'b00000000,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00000000,8'b00000000},
        '{8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b00000000,8'b00000000,8'b11000000,8'b11000000},
        '{8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000000,8'b00000000,8'b00000011,8'b00000011},
        '{8'b11111100,8'b11000000,8'b11111100,8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11000000},
        '{8'b00111111,8'b00000011,8'b00111111,8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00000011},
        '{8'b11000000,8'b11000000,8'b11000000,8'b11000000,8'b11111100,8'b11000000,8'b11111100,8'b11000000},
        '{8'b00000011,8'b00000011,8'b00000011,8'b00000011,8'b00111111,8'b00000011,8'b00111111,8'b00000011},
        '{8'b11000000,8'b11000000,8'b11000000,8'b00000000,8'b11000000,8'b11000000,8'b11000000,8'b00000000},
        '{8'b00000011,8'b00000011,8'b00000011,8'b00000000,8'b00000011,8'b00000011,8'b00000011,8'b00000000},
        '{8'b00111100,8'b00111100,8'b11111111,8'b11111111,8'b11111111,8'b11111111,8'b00111100,8'b00111100},
        '{8'b00000000,8'b00000000,8'b00111100,8'b00111100,8'b11111111,8'b11111111,8'b00000000,8'b00000000},
        '{8'b00000000,8'b11111111,8'b11111111,8'b00000000,8'b00000000,8'b11111111,8'b11111111,8'b00000000},
        '{8'b00011000,8'b00011000,8'b00011000,8'b00011000,8'b00011000,8'b00011000,8'b00011000,8'b00011000},
        '{8'b00011000,8'b00011000,8'b00011000,8'b11111111,8'b00011000,8'b00011000,8'b00011000,8'b00011000},
        '{8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100,8'b00111100},
        '{8'b00000000,8'b00111100,8'b01111110,8'b01111110,8'b01111110,8'b01111110,8'b00111100,8'b00000000},
        '{8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000}
    };

    // VGA Output
    always @(*) begin
        VGA_R = 0;
        VGA_G = 0;
        VGA_B = 0;

        if (tile_bitmaps[tile_id][ty][7 - tx]) begin
            VGA_B = 8'hFF;
        end
    end

    // Tile initialization
    initial begin
        integer i;
        for (i = 0; i < 4800; i = i + 1) begin
            tiles[i] = 0; // Default to background
        end

        // ====== Your tile assignment here ======
        tiles[35] = 23;
        tiles[3765] = 12;
        tiles[4500] = 8;
        tiles[1800] = 15;
        tiles[2500] = 5;
        // You can continue your 2000 lines here
        // ========================================
    end

endmodule
