2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h2 2'h2 2'h2 2'h2 2'h2 2'h1 2'h2 2'h2 2'h2 2'h2 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h0 2'h0 2'h0
2'h0 2'h1 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h2 2'h2 2'h3 2'h3 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h0 2'h1 2'h1 2'h1 2'h0 2'h0 2'h1 2'h1 2'h1 2'h0 2'h1 2'h1 2'h0
2'h0 2'h1 2'h0 2'h0 2'h0 2'h1 2'h1 2'h0 2'h0 2'h1 2'h1 2'h0 2'h0 2'h0 2'h1 2'h0
2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0
