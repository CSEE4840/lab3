00000000
00003C00
00FFFF00
03FFFFC0
10E4791C
11CB2E74
11D33B74
75D33B7E
787479DE
7FFFFFFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
6E1C3B1A
43198642
00000000
