// left
0000
07C0
1FF0
3FF8
3FF8
0FFC
01FC
00FC
01FC
1FFC
3FF8
3FF8
1FF0
07C0
0000
0000


// up
0000
0000
1830
3878
3C78
7C7C
7C7C
7EFC
7FFC
7FFC
3FF8
3FF0
1FC0
07C0
0000
0000

// down
0000
0000
07C0
1FE0
3FF0
3FF8
7FFC
7FFC
7EFC
7C7C
7C7C
3C78
3878
1830
0000
0000

// right
0000
03E0
0FF8
1FFC
1FFC
3F80
3F00
3F80
3FF0
3FF8
1FFC
0FFC
07F8
03E0
0000
0000

//eat
0000  
07E0  
1FF0  
3FF8  
3FF8  
7FFC  
7FFC  
7FFC  
7FFC  
7FFC  
3FF8  
3FF8  
1FF0  
07E0  
0000  
0000  

