0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0002
0001
0000
0001
0001
0001
0000
0001
0002
0001
0000
FFFF
FFFF
0001
0000
0000
0001
0000
0001
0001
0000
0001
0001
0002
0001
0002
0002
0000
0000
0000
FFFF
0000
0001
0003
0002
0002
0003
0002
0000
0001
0003
0004
0003
FFFF
0002
0004
0000
0003
0008
0006
0006
0005
0002
FFFF
FFFE
0001
FFFF
FFFF
FFFB
FFF4
FFF8
FFFB
FFFA
FFFC
FFFB
FFFB
FFFB
0000
0002
0008
0010
0006
0004
000E
0008
0004
0004
0009
000C
0001
FFFA
FFFB
0003
0006
0004
0008
0006
0004
FFFF
FFFD
0003
0002
000C
0013
0005
0001
0006
0004
0000
0003
0005
FFFD
FFFF
FFFB
FFFE
000A
FFF7
FFF4
FFFC
0008
001F
000B
0001
0006
0002
0017
0009
0005
0027
0009
FFE4
FFF0
FFF6
FFF0
FFFA
FFEB
FFD2
FFF0
FFE5
FFD4
000A
FFFF
FFFB
001F
0009
001A
0026
000E
001E
001B
0011
FFF9
FFE0
FFFB
FFF6
FFF4
0016
0011
000C
0016
0013
0007
FFF7
FFF7
FFFB
FFEF
FFD5
FFD6
FFF6
FFF2
FFE9
FFF0
FFDC
0008
0049
0024
0000
0001
FFF6
0004
0001
FFDE
FFD4
FFE5
FFEE
FFDA
FFD7
FFE7
FFFB
000C
FFF7
000E
0021
FFF5
000C
FFF4
FFBB
FFD3
FFCC
FFE9
FFFD
FFEF
0028
0013
0015
0049
0021
0044
004F
0010
002D
001F
FFE2
FFE5
FFFA
FFF5
FFF4
FFDA
FF8D
FFBD
FFF9
FFC5
FFFE
0012
FFE8
000A
FFDC
FFED
0032
0018
0014
FFDA
FFCC
0011
FFEB
FFCE
FFD0
FFCE
FFFA
FFF7
FFE6
FFFB
FFFC
FFD8
FFD4
000C
0006
FFED
0004
FFE1
FFB9
FFC6
FFEC
0015
000B
000D
0021
0000
FFE2
FFDF
FFFA
0013
FFF0
FFEF
0026
0017
FFEA
FFF4
0015
0036
0049
0048
002F
0005
0015
0052
006D
0056
001F
0010
002C
0042
0021
FFD9
FFEC
FFF4
FFCF
0010
FFF6
FFB5
000D
001B
000D
0035
0015
000B
001B
0014
0009
FFE2
FFEA
0022
0031
0028
002E
0018
000C
002D
000E
FFE7
FFE2
FFDE
0016
0000
FFCD
FFF1
FFFC
0039
0035
000A
0050
000A
FFEC
0020
FF9C
FF9B
FFF4
FFF2
0027
0017
FFD1
FFF0
0006
FFAE
FFBF
0023
FFD6
FFD3
0018
0013
0071
0038
FFDE
0005
FFDF
0021
0018
FFD1
0021
000B
001B
0008
FFBC
FFEE
FFAE
FFDF
0014
FFCE
0046
001A
FFCC
FFFE
FFCD
0001
FFD1
FFBD
0024
FFDC
FFDA
FFE4
FFE1
FFDE
FFAE
FFE7
FFA8
FFF0
002D
FFB0
003C
FFEB
002E
004A
FF60
014B
FF0C
00E4
11CA
19A5
148A
1376
1159
0EDC
0E5C
0C07
0B44
0A68
08B9
07E8
068C
05BC
0486
037F
02FF
01A3
013D
005C
FF3E
FF1C
FE06
FD8C
FD16
FC20
FBF3
FAF3
FA7A
FA56
F95B
F93C
F8F0
F887
F830
F775
F7A0
F77C
F712
F6E7
F68B
F6AB
F623
F5FB
F682
F649
F695
F607
F5C7
F68A
F5C8
F64F
F62A
F594
F6D5
F513
F72B
F5E4
E3B9
D9E3
DF8E
E162
E38D
E67D
E75B
EA27
EB25
EC5E
EE46
EF0B
F15C
F294
F3D8
F592
F5CE
F77C
F8C2
F975
FAFE
FBCF
FD14
FE04
FEDE
0012
00AB
0203
02B8
0340
0474
04C0
0589
0605
0655
0736
077C
0874
091D
0988
0A2B
09E5
0AD7
0B61
0B1E
0B93
0B73
0C71
0CB3
0C8A
0DB7
0D02
0D96
0DAA
0CFC
0F0E
0C39
118C
24DE
2A04
242A
234A
209C
1E7E
1D81
1B1F
1A9F
190C
178C
16AB
148A
13CB
129A
112B
1083
0EDB
0DDF
0CDB
0BAC
0B14
09E7
0912
07EF
06FE
0696
0562
04D0
040B
0324
02C4
019D
0127
0095
0000
0010
FEE1
FE4B
FDD5
FD43
FD53
FC11
FC07
FC43
FB58
FB4F
FA67
FA65
FA6A
F9BF
FA64
F915
F961
F94A
F7C5
FAF7
F163
DE9E
DD98
E283
E342
E676
E7B3
E8F8
EA8F
EAFD
ED0D
EDD1
EF12
F0FE
F162
F2E8
F3C1
F490
F64B
F6A6
F7D1
F921
F986
FA82
FB43
FC13
FCD8
FD7D
FE30
FEB5
FFD7
0055
0079
0129
0171
0221
0298
0300
03C1
03B7
0465
04A7
048B
0591
0573
0587
05D3
05D0
06A0
0633
0690
06E6
0672
079B
0678
0760
07B3
04F3
1292
22F6
2036
1CD6
1BFB
181D
1770
1592
1405
136F
10EF
1067
0F19
0D6B
0D02
0B2B
0A3A
0901
0750
06D0
0566
0442
0373
0292
0209
00D6
0041
FF81
FE7D
FE44
FD3E
FC79
FC1B
FB5E
FABC
F9D2
F97A
F90A
F866
F85B
F7B0
F751
F728
F6BA
F687
F5F8
F602
F57A
F508
F582
F474
F4B6
F4B3
F3FB
F58C
F36C
F47D
F563
E438
D75F
DC50
DE88
E00B
E364
E3B0
E5D4
E738
E849
EA96
EB2F
EC89
EDCA
EEA1
F033
F12D
F2A0
F3A7
F47D
F5C8
F686
F7D7
F89C
F93F
FAA0
FB47
FC0D
FCC8
FD5A
FE13
FEBA
FF89
FFC5
009D
0164
017B
023F
0233
02EA
040C
03D6
0446
0495
057B
05CC
059C
06C1
05C7
0791
0528
F80B
F599
F985
F8CA
FD10
FC2C
FF06
11C3
197A
1559
151D
13BB
1294
1287
1191
11C9
1134
101E
0F71
0ED8
0EB8
0E1E
0D8C
0CDB
0C3A
0C2F
0B6E
0B19
0AF3
0A0B
09B2
0936
08AE
086E
0820
07CD
06D3
06AE
06AC
05A4
058B
0565
0504
049B
0416
0476
03B0
0340
0360
028B
02A9
0162
013F
01BD
000A
016D
FF24
01D0
11AB
148E
1011
1065
0BC4
0D30
064F
F095
EC4D
F0A6
EFCF
F236
F2AF
F2D0
F3B1
F36A
F496
F49C
F543
F5E1
F562
F68D
F6C2
F716
F7AC
F781
F84A
F867
F8DD
F93D
F929
FA13
F9D1
FA5E
FB2F
FAD3
FB89
FB46
FBBB
FC9E
FBC6
FC59
FC91
FCB8
FD8D
FD45
FDE4
FDCC
FE17
FEF7
FE6F
FF71
FEC5
FE8D
FFD5
FE96
00F8
FBF3
EF0C
EF34
F17F
F205
F5C0
F3A3
FDB5
0FB3
0FC8
0CDC
0D6B
0AE7
0B1E
0A6E
0978
09DC
088D
088F
0853
0784
0768
06A9
06A5
0632
05AA
059F
04CD
04C0
0456
03B3
03A3
030D
0301
02AF
0265
0290
0235
0219
0157
0135
0182
00E8
013B
00B6
008C
00A6
FF44
FFEF
FFAF
FF04
FFB7
FEB3
FF45
FE96
FE8C
FF86
FC8A
0673
13B5
10B7
0F6E
0DB1
0AED
0C88
FC39
EB8B
EEB0
F062
F0AE
F2FA
F295
F409
F4A1
F4C0
F569
F5A1
F719
F715
F768
F850
F831
F92F
F933
F9C1
FB02
FAAA
FB80
FBDB
FBF4
FD1B
FD1E
FD6C
FD9E
FDF7
FEAE
FE61
FF20
FF58
FF0F
FFF5
FFE8
004E
00DE
00F6
0177
018B
0220
0210
0240
0291
0216
03BB
026E
028A
0487
F92D
F0FB
F4EE
F528
F839
F8B2
F8F8
0AA2
1575
1179
1140
1001
0EDC
0F3E
0D5D
0D98
0D19
0C26
0C69
0B1F
0ACD
0AB6
0A0D
09AD
0924
0946
08AD
0839
0838
0764
075C
0705
066D
064B
05E8
05F6
0542
04F6
0500
03FB
042C
042A
03C3
03C1
0325
032F
0286
026A
02A0
0150
01F9
0190
012F
022B
004F
0138
FFF5
00F9
0FF9
15BA
1102
10E3
0D0A
0E2F
09F9
F45E
ECC7
F176
F113
F35A
F3FA
F39F
F55B
F4D7
F5B5
F669
F687
F798
F769
F7ED
F840
F8D0
F9D2
F957
FA48
FAF9
FAEE
FBB3
FB6F
FC0D
FC9D
FC4A
FCD7
FCF7
FD73
FD96
FD73
FE2E
FE37
FEC1
FED6
FE6F
FF19
FF48
FFDA
FFEC
000D
00A8
FFDE
00E5
00E9
005D
019B
004A
026D
FF08
F18B
F05F
F395
F362
F769
F54F
FCA2
0FCF
11FB
0E31
0F05
0C9B
0C79
0C0B
0AB5
0B23
09FC
09E3
09B4
0892
0828
0752
0765
06CC
0609
064C
055F
052F
0506
047E
046A
0368
0391
0353
024D
027D
0196
016D
01C6
0128
0131
007A
007B
00A8
FFB7
FF8F
FF15
FF35
FEB9
FE0C
FED5
FDF3
FE7B
FE2E
FD1E
FE8A
FBAC
02B9
117F
1032
0DAC
0CE0
08E4
0B41
FE30
EA66
EB6C
EE7B
EE6F
F0EC
F063
F18D
F25E
F20B
F32F
F36A
F440
F47E
F4D6
F591
F543
F663
F674
F65B
F772
F70E
F7DA
F88D
F884
F99E
F9A7
FA05
FA7E
FA6E
FAE8
FAE0
FB6D
FBAB
FBAF
FC65
FC41
FCFB
FD5A
FCFB
FDA9
FDE9
FECD
FE8A
FE0F
FF06
FE18
FF40
FF54
FE71
00EB
F7AD
ED15
F090
F184
F32F
F544
F465
03EA
11A3
0DB5
0CA5
0CA8
0AB1
0B2E
09C8
09A3
09C4
08BF
089E
0799
0758
06A3
05BD
062E
055C
0539
0518
043F
046A
03E8
039A
0305
0268
02BE
0209
023B
0255
0158
013A
008F
00C9
00DB
000C
007C
FFCF
FF85
FFD1
FF60
FF8C
FEA9
FE96
FE53
FDB4
FE8D
FD0B
FE08
FDC3
FCEF
0AAE
1353
0E92
0E40
0AE3
0A6B
08F1
F4C1
E9E0
EEB5
EE92
F03D
F1F3
F166
F379
F387
F40B
F4CA
F454
F581
F5CE
F64B
F6E1
F6E0
F811
F868
F8FA
F980
F96F
FA78
FA66
FAB2
FB52
FB0C
FC45
FC6C
FC26
FD4A
FD35
FD3C
FDB9
FDEB
FE2A
FE5F
FEF5
FF3A
FFCA
FFE8
FFDE
0077
FFBB
008C
0129
008D
0209
0106
026F
0140
F435
F01F
F403
F426
F7E5
F6A3
FB77
0E9E
13E2
0FC3
0FFF
0DB1
0D35
0D5A
0BF1
0BF8
0B1F
0B2A
0AE9
09C2
09ED
095B
08F4
0899
07E8
0850
08DC
0924
0841
0790
077D
0649
063A
062C
0546
0559
04C0
0408
03C2
0369
0332
02B8
0329
030A
01F0
0201
021D
01C8
00E7
00A4
0111
007D
0088
FF7F
FF25
0073
FE11
03B2
11EE
1403
0FAC
0EAE
0C0C
0AF3
08FE
04F3
0475
03C2
02B9
02CD
0177
00FB
0069
FF32
FEDE
FDDF
FD92
FD40
FC71
FC91
FBAF
FB64
FB14
FA6D
FB4C
F9A5
F9A7
FA98
F7FE
FAA3
F54C
E24D
DD30
E264
E311
E5A8
E7AD
E8A3
EACE
EB22
EC8B
EE93
EF7E
F0EB
F209
F325
F429
F4BB
F5F8
F6FA
F797
F956
F9E3
FA73
FCED
F658
EB32
ECCE
F145
F1C6
F544
F6EA
F7A4
F974
FA51
FC3F
FCF8
FE1E
000D
009A
0290
0370
044E
061F
0615
0767
0840
0889
0A28
0A80
0B81
0BED
0C46
0DBC
0D5C
0E58
0EAA
0E4D
0FD1
0F1E
100B
1067
0F9D
11F5
0F55
149C
2634
2A28
2531
242D
21CC
202C
1F4A
1DF3
1D30
1B83
19CE
18EB
180E
15FE
158A
1431
1255
1CC0
270D
2302
1F61
1D9E
1A03
184A
159F
13F2
124F
0FBA
0EB9
0CBA
0B1C
09BB
07F3
06FD
050E
0419
02FB
0127
004B
FE80
FDDE
FCBF
FB08
FB4C
F9D0
F8C6
F811
F66A
F6D7
F5E7
F4F9
F4B8
F3A1
F3C9
F28B
F22A
F21D
F0D9
F15D
EFD0
F02E
F06F
EEAF
F1B1
E6BE
D47A
D54E
D935
DA2C
DD74
DDB5
DFEB
E09F
E24C
E3BE
D93E
D3F5
D94D
DB26
DDB2
E0D6
E274
E513
E6B4
E880
EA19
EB7E
EDA2
EF74
F16D
F29E
F41B
F618
F70D
F8D4
FA4B
FB24
FC73
FD46
FEAD
FFCD
008A
01DC
02F8
0433
0489
0510
0646
067E
079D
083D
085A
09AD
09A4
09EA
0AB5
0AE6
0BC7
0BDD
0C15
0C49
0C88
0D5D
0CC4
0D6D
0D33
0D2B
0EBA
0BE5
1560
269A
2368
236B
319D
3281
2D0B
2AF5
272A
24CF
224D
1F61
1D89
1B61
19A4
17A7
1587
1343
1110
0FC0
0DFC
0C1A
0A9A
0933
079D
05BC
0493
0333
016D
002B
FED1
FDAB
FC96
FB7A
FA6D
F94C
F874
F79A
F6EF
F618
F529
F4D3
F416
F373
F314
F286
F244
F189
F0E5
F093
F01F
F00A
EFBB
EF11
EEBB
EF13
EEBD
EE66
EEDA
EE1F
EF7C
EA2B
DA5F
D9B7
DEE8
D09E
C774
CD14
CFFD
D302
D6A3
D846
DAFE
DD44
DFBC
E28F
E45E
E64F
E8AF
EAE5
ECAC
EEE6
F0FE
F24B
F3C8
F538
F707
F89B
F999
FB85
FCB9
FDCC
FFD2
0066
0116
027C
034C
047A
053A
062B
0778
07CB
0888
095B
0A13
0AD7
0AFB
0BEF
0C5C
0C72
0D76
0D68
0DC7
0E60
0EA8
0F92
0F38
0F94
1021
0FB7
1013
0F87
1017
1036
0FBE
10F4
0F4D
105C
1083
0F2D
1E02
29C2
2512
2371
21CF
1F10
1E68
1BD9
1B17
1947
17E2
1714
153C
154E
1195
164D
2364
229D
1E15
1CCA
1934
17D0
153B
130F
119E
0ED1
0DFA
0BB5
09E0
08ED
0661
0573
03E9
025D
0170
FF9E
FED6
FDA1
FC97
FB56
F9F1
F9B2
F812
F751
F6DF
F5B2
F5F4
F501
F49C
F43A
F2EF
F330
F225
F180
F118
F033
F096
EF72
EFA8
EF6F
EECB
F028
EDBC
EFF2
ECD1
D908
D270
D811
D820
DB4A
DD89
DE82
E122
E182
E37D
E4B9
E650
E7CE
E7C4
EB81
E682
DBBB
DCFE
E0BA
E29B
E609
E78A
E9D2
EC19
EDA7
EF94
F115
F356
F4D3
F67C
F85E
F902
FABA
FC1C
FD7B
FF36
FFE4
0178
0278
031E
048C
055A
0686
0747
082A
08EA
091D
0ACD
0B3B
0B7D
0C7D
0CA4
0DBF
0DA3
0E3C
0F4F
0E66
0FCD
0FD1
0FB8
10A4
0F79
11AE
0FFD
12CA
2479
2A55
2563
24D6
21D5
2097
1FD3
1DCF
1D46
1B00
1A5D
18BE
17A3
16E4
13FA
1E16
28D4
2487
2184
1F6D
1BD5
1AA0
17C3
162D
1458
11E2
10ED
0EB7
0D4A
0B6B
09B3
0919
06DE
05C7
0466
0292
020A
0058
FF7E
FE65
FCD3
FC92
FB3D
FA58
F9B4
F8FB
F87E
F6FD
F6D3
F648
F566
F56A
F41E
F3F9
F364
F2E4
F371
F1D5
F22B
F1AA
F0DB
F21C
EFC1
F226
EE37
DA60
D427
D9B3
DA99
DDA8
DF51
E07D
E2D8
E351
E537
E627
E797
E8AB
E9EB
ECCB
E485
DBF5
E002
E260
E3F8
E779
E8DF
EBA7
ED70
EF3C
F19F
F26F
F453
F5E5
F78A
F950
FA1D
FBFB
FD26
FE12
FF96
00C2
0257
02EE
03D5
0554
0605
070C
07BE
0845
08DE
09A9
0A72
0AAF
0C08
0C8C
0CBB
0DBC
0D94
0E95
0EC1
0E9A
0F9A
0ED6
0FF5
0FDB
0FC7
11AE
0E7B
1701
27FB
2808
241E
2377
2039
1F90
1E07
1C71
1B7D
19E8
192D
16FB
170F
14CA
1482
216E
275E
21CA
1F9F
1CB9
1A0E
18AC
15F7
1460
11FB
0FFC
0E87
0C88
0B3A
091E
07CB
0692
04AB
03CB
0231
0105
FFC6
FE19
FD9A
FC1B
FAF8
FA27
F8C6
F84A
F72A
F6B4
F60E
F4A8
F4EE
F40F
F31D
F2A6
F1CD
F202
F0D8
F09B
F0A3
EF61
F001
EEF4
EF43
EF58
EDB6
F0FD
E6CC
D3E5
D3D2
D844
D8E1
DC35
DD57
DF5E
E0B9
E1AD
E3DB
E497
E70C
E779
E99A
EA5D
DEDA
DA20
DF93
E135
E3F9
E61F
E7C8
EAEF
EBFE
EE4D
F03B
F1A9
F3DC
F4BC
F6C5
F814
F91E
FB45
FC30
FDB3
FEE2
FFE4
0179
0214
0313
03EB
04F9
05D0
05FC
0771
0833
08DD
099F
09F4
0AFD
0B12
0BDE
0C4B
0C59
0E09
0D8E
0E00
0EA8
0E56
0FB9
0E29
0FBB
1031
0DAA
1BE9
28F0
2510
230B
2165
1EF1
1E5F
1C6A
1C1F
1A42
18E4
1818
161C
165D
1292
1668
244E
24D9
1FB9
1E5A
1AE2
194E
171F
14AD
138C
10F1
0FBC
0DCA
0B82
0A6C
0864
077E
060C
0421
0300
014E
00CC
FF83
FDCC
FD29
FBA8
FAE8
F9E6
F8C7
F853
F704
F6D4
F641
F51C
F4D7
F423
F411
F319
F24A
F24D
F14A
F18D
F095
F031
F0AE
EF15
F09C
EF60
EEFF
F0F4
E112
D2A3
D6EA
D922
DAD3
DE06
DE7B
E0D9
E185
E2FF
E522
E61B
E7EA
E810
EB78
E8AE
DCF7
DCBB
E16A
E2CD
E66C
E7E7
E9C7
EC2F
ED56
EFDC
F121
F2FB
F4DB
F5C8
F804
F92A
FAD5
FCCA
FDA1
FF30
FFDE
00F5
0256
0332
04B3
0529
0636
07B3
0813
08DC
098F
0A47
0ABC
0B4D
0BFE
0C40
0DA2
0DCA
0DCA
0ED1
0ED1
0FB9
0F74
0FBE
10C2
0FCD
11EA
0FD6
115D
22AB
29F8
254C
24BD
21D6
2010
1F1D
1CE3
1D13
1A98
1979
1897
169A
1732
135E
17E1
25DD
2616
2106
1F9B
1BEB
19EE
181F
15AF
13F1
119F
106B
0E99
0CB3
0B9B
097E
0806
06E1
056F
03EB
0310
031E
0163
FFE5
FF58
FDD7
FD2D
FBFA
FAA1
FA3D
F903
F82F
F765
F684
F5D1
F4D9
F4B4
F3D9
F33C
F34F
F244
F1DA
F133
F0B5
F0A8
EFE8
F04E
EFA6
EF54
EF5C
EC2E
EB44
EC12
EBDA
ECBB
ECD4
ED3E
ED12
ED04
EE2E
ED9A
EEDB
EEB5
EE75
F0EC
E6D2
DA9E
DD2F
E02F
E121
E402
E4F5
E713
E8D6
E9A7
EBB7
EC84
EDCC
EF79
F034
F1E2
F2C9
F411
F5D5
F58A
F790
F87E
F851
FC20
F3EF
E513
E658
EB36
EC59
F014
F1B3
F3FB
F688
F75D
F9C5
FB2E
FC8D
FE87
FFE1
01A6
02B7
0420
057B
068B
0836
08F4
09BE
0ADD
0BF9
0CF8
0CFF
0DCD
0EE1
0F48
1001
1091
1102
11DA
1224
123A
1341
132D
13A0
1420
1319
1BA1
265F
249D
22AE
2291
2004
1F78
1E1E
1D8A
1CD6
1B34
1B26
1950
18A9
1812
168B
169F
1532
1482
13B1
12BC
1272
10BB
1125
0F73
0F22
0F28
0B61
190C
28A8
2402
209E
1EB1
1A55
194D
1650
14D5
1308
1024
0F24
0CD4
0B41
09BE
081C
06E0
04F2
040D
023B
00F8
FFFA
FE2E
FD6C
FB9D
FB50
FABB
F904
F8FF
F6DE
F64B
F5F4
F43B
F525
F2C4
F344
F2A6
E43F
DBB9
DF61
E087
E153
E320
E394
E45E
E513
E5B7
E6B5
E741
E80D
E8EF
E91F
EA3A
EB55
EBE4
ECBA
ECED
EDDD
EE7B
EF09
F056
F036
F13A
F12F
F18F
F38C
F18B
F46D
F2D5
E1D8
DBFF
E1C8
E300
E5B5
E866
E9A5
EBCD
ED50
EF71
F0F5
F23A
F3D3
F4E6
F622
F742
F8C9
FA15
FB25
FC9A
FD71
FE30
FF62
006A
010D
0224
030C
038B
0465
047D
0600
05D1
06E0
12F3
1A58
16BF
1671
15BB
140D
1415
12FE
1307
1226
1187
117E
102B
0FF8
0EEF
0EAD
0EA9
0D08
0D0A
0C30
0B88
0B45
0A4C
0A98
097A
092F
090E
0818
08C0
0739
0748
06CC
052B
0717
036D
094F
1CC0
1FC8
1A39
194C
15A7
1382
11D4
0FAD
0EAB
0C7F
0B19
0974
07B1
06CA
0572
0423
0280
014E
0015
FF53
FEBC
FCB6
FC00
FAD9
FA26
FA21
F7CD
F97A
F4F4
E559
E13A
E52B
E4DA
E698
E7DA
E7CD
E930
E96B
EA0A
EADC
EB23
EC08
EC92
ED42
EE0F
EE68
EF77
F056
F06F
F133
F1E4
F224
F2E4
F3AA
F430
F48C
F52F
F5C1
F654
F7A0
F766
F7B2
F8D3
F86A
FA78
FA98
FA82
FCBA
F051
E2B7
E665
E961
EA8E
EE53
EEF4
F11D
F2A3
F383
F5C2
F691
F8A7
F9BE
FA69
FC91
FD11
FE58
FFCD
00A7
01FB
0246
0338
0466
0579
0607
05C8
0718
078A
07DB
0931
0924
09DF
0A8F
0AAF
0B78
0BA8
0C58
0CA9
0CD6
0D9F
0D97
0E09
0E82
0EA9
0EF5
0ED9
0F26
0F17
0F3A
0F71
0F0C
0F96
0F9A
0F65
0FB5
0F33
0F25
0F12
0EBE
0ED8
0EA5
0EE9
0E5E
0DD1
1538
1FBB
1CA4
19FA
2A19
342C
2E5E
2B17
282E
242A
2241
1F32
1D1B
1ACE
185E
16E3
141B
1245
104A
0DC3
0C62
0A62
08BE
0704
051A
044F
0301
0175
0033
FF14
FDE1
FC0B
FAD2
F9DE
F8AD
F7B4
F6D2
F635
F56B
F45B
F348
F28A
F249
F1CA
F12D
F072
EFF2
EF97
EF09
EEFD
EE6B
EDAE
ED96
ED51
ED87
ED79
ED03
ECD5
ECAC
ED57
ED12
EC3E
ECBE
EC91
EC86
ED01
EC63
EDA5
ED61
E1CF
D6FC
DCC0
DD2A
CDCD
C8E4
CEBC
D1A4
D51B
D82B
DA80
DD9D
DFC2
E257
E4A0
E6B5
E924
EB2B
ED79
EF2F
F0FE
F323
F4B8
F68A
F7F3
F98E
FB77
FD06
FE87
FF58
00F7
02C3
039B
0529
0621
0703
0860
08CF
09CC
0AEC
0BC1
0C99
0CC9
0DB7
0ED2
0F04
0F4C
1005
10FE
113F
116D
1202
120E
1285
1308
1304
1368
13A8
139A
137C
1396
1422
1423
13D3
13A0
13DB
1456
1306
16AE
2369
2641
1F04
28C6
38D5
379F
3236
300A
2BE3
2932
26B5
23EE
2212
1F30
1D04
1B25
18B2
16C9
148C
1267
10B2
0EF3
0D17
0B54
09EB
084A
06C7
052A
0391
0275
00D7
0004
FF35
FD52
FC6D
FB1C
FA0C
F9EC
F836
F738
F704
F5E2
F55D
F48D
F3B6
F388
F2DD
F229
F1A6
F153
F118
F07C
EFDF
EF9C
EFB3
EF92
EF2A
EEDD
EECA
EEE7
EE94
EE88
EEA4
EE17
EE4D
EE09
EDF1
EFAC
E8E9
DA72
D9E1
DFEF
D4AA
C8B2
CC92
D146
D360
D6FB
D95D
DC3F
DEBC
E0CB
E384
E52D
E791
E9F0
EB78
EDB7
EF62
F106
F2E9
F492
F678
F7D1
F975
FB23
FC3E
FDD9
FF3C
0078
01CC
027E
035A
04B7
05C9
064B
0709
082C
091E
09C8
0A13
0AB6
0BF4
0CB4
0D0D
0D8A
0DF0
0E75
0F5C
0F8D
0F40
0FB5
0FFF
100A
104C
1078
10C1
1097
108F
10D7
10A1
10E0
10EC
1088
10FC
1068
10EB
1A80
23D4
1E66
1EFE
30F4
3758
308E
2DF3
2A9B
26E0
24F0
21CB
1FAA
1D3A
1A96
18BE
168E
14B0
125E
1054
0E92
0C78
0AF0
0914
0784
05CE
03AD
02CE
015E
FF91
FE94
FDA1
FC98
FAF6
F9BA
F8CB
F77B
F6FB
F65F
F540
F473
F3D1
F322
F24A
F1D4
F147
F06C
F002
EFB3
EF3E
EEC2
EE71
EE1B
EDA9
ED89
ED5C
ED32
ECE5
ECB5
ECE9
EC85
EC70
ECB1
EC2E
EC6B
ECAC
EC0B
ED89
EBB6
DE39
D5F1
DD7C
D9FE
CA34
C8A1
CE5E
D07E
D427
D74D
D9E4
DCCC
DEA1
E0DA
E316
E557
E7C6
E9F4
EC16
EDAA
EF75
F176
F319
F4DB
F691
F851
FA1A
FB67
FCBC
FE8C
FFAC
0074
024C
0360
03CA
0552
0687
0753
081F
08AB
099D
0A98
0B67
0C10
0C9A
0D21
0D93
0E3B
0E82
0F0C
1007
1029
1059
10D3
10CE
10CD
113A
119D
1189
11A8
11D0
11EC
11E1
11B7
120B
11E1
124A
1167
13C3
2111
2470
1DA7
2ADD
3932
34E7
30C8
2DD3
29F7
284E
24B7
225A
207E
1D7D
1B9A
196E
1741
14F9
12FC
1140
0F02
0D8E
0B8E
09D2
08BC
06B6
057E
03F0
0227
015F
003A
FF44
FDE1
FC86
FBE4
FAA6
F9B8
F8C5
F7DF
F745
F62C
F596
F4BD
F3D0
F367
F2A9
F24C
F193
F123
F152
F07E
F036
F001
EF4A
EF3E
EF28
EF6C
EF1D
EE5E
EEEA
EEEF
EE9F
EEB1
EE77
EED3
EE79
EEC8
EF98
E69A
D9BB
DC66
E039
D281
C8E9
CDE6
D212
D4DD
D874
DA93
DD68
DFD5
E220
E4C2
E692
E8FF
EB04
ECBB
EF25
F0C5
F264
F481
F664
F7D4
F944
FB47
FCB9
FDF6
FF95
00F4
024E
032C
0457
059C
0636
0789
087F
092D
0A55
0B0D
0C0B
0CA6
0D2F
0DD9
0E26
0F77
0FCF
0FE3
1088
104E
1166
1187
1187
1316
13DA
15E3
1447
15F4
234E
2884
24C0
23E7
21D8
2071
1F02
1E2F
1CFE
1B1C
25F4
2F34
29AA
27B9
2875
2623
2418
2081
1E9C
1CF3
1A1C
180A
15AC
144B
123C
1060
0F5A
0CC3
0B41
098F
076D
069F
04C5
0388
02B2
0130
002E
FEAA
FDA7
FCCB
FB7D
FB05
FA27
F910
F85A
F783
F6B7
F608
F595
F4C7
F408
F38F
F2FE
F2F7
F26C
F1A2
F171
F0DD
F0F4
F0E9
F00A
F022
F026
F03F
F01F
EF2F
EFED
EFA5
EF63
F05A
EE84
F0EA
ED3A
D9DF
D469
DAEA
DA54
DF8C
DE54
D217
D202
D67A
D873
DC6F
DE7E
E103
E3B4
E577
E7F0
EA2A
EC6F
EE09
F00D
F229
F39F
F5EE
F75D
F8FB
FAB0
FBA8
FD58
FE15
FF75
0152
01B9
02DD
044A
05A4
06BE
07C1
08FA
092F
09FB
0AA6
0B21
0C25
0C47
0D44
0DD2
0E06
0F2A
0F0F
0FC0
1065
10A6
1179
112E
11A4
11BD
11AD
1224
117D
120B
11E4
11E9
126A
117E
1282
11FB
11C6
128A
112F
1294
113F
112E
12AB
0E94
167F
1FA1
22CA
3334
395F
310C
2EE7
2AA6
275A
2600
21FD
203F
1D59
1AB5
1902
1678
14CF
11F3
1007
0E86
0C35
0AC9
0864
06D2
057D
0386
0246
005D
FF11
FDAB
FC24
FB98
FA0A
F8DE
F7FE
F6CE
F5D5
F490
F421
F332
F1F1
F166
F08E
F062
EFCE
EEDD
EE75
EDA1
ED7D
ED28
EC77
EC6B
EC38
EBDF
EB57
EB45
EB78
EB64
EAF1
EA4D
EB0C
EB19
EACB
EB0B
EA56
EB54
EA8D
EAB3
EBAB
DF2D
D55E
DA09
DB21
DCF6
E018
DF98
E2D9
E2D1
E4A9
E738
D952
CF43
D484
D7D1
DA70
DE36
E05E
E2E7
E4BF
E719
E95C
EAEF
ED25
EED4
F0F7
F314
F4B5
F6A3
F7D3
F993
FB5F
FC82
FE5F
FFB7
00D8
020B
031A
04C3
0599
0699
07F5
0834
0906
0A0C
0ABC
0BDA
0CE3
0DB1
0DC0
0E27
0F17
0F48
0FDA
1039
1061
10F4
1112
11C3
1203
11C2
1253
1234
12BF
12B3
11FA
139B
1229
1364
1F48
2548
216F
205C
1EF6
1CB4
1CA2
1AFE
1A3E
19CF
17EF
17BE
160A
14B1
1501
12BD
1311
1135
0EF1
1DD2
2B2A
262C
2238
2063
1C31
1AF1
1823
15B7
14AF
1218
10E6
0EED
0C96
0B45
0941
081E
061F
0413
0314
012B
0080
FF77
FDA9
FCA3
FB18
FAF2
F9C2
F7EC
F817
F648
F5DE
F5BC
F392
F558
EF32
E03C
DD5A
E0FD
E0CF
E2BF
E448
E41E
E524
E5BA
E67B
E742
E813
E925
E987
EB44
EC8F
EC54
ED5E
EDD4
EE53
EF81
EF85
F026
F0D6
F14F
F208
F269
F33D
F343
F3E4
F4D7
F4BB
F605
F626
F687
F78F
F6F0
F8E7
F84C
F8C3
FB84
EE4D
E14B
E52F
E816
E992
ECC1
EDA9
F01B
F19B
F2A5
F4AF
F5C3
F775
F8CE
F9EA
FB18
FC09
FDA3
FEF1
003E
0139
01CF
02B0
03C5
04F1
0524
063D
06CB
0706
08DE
07BB
0D33
1991
1AB2
1828
1899
1679
1647
15CD
14F3
14DB
12ED
12D6
1249
1129
11BB
10EB
1065
0FEF
0F71
0F1D
0E06
0E53
0D9C
0CAD
0D02
0C33
0C1F
0BD0
0BA6
0B9F
0A54
0ABF
09F9
08E0
0934
0812
0821
0791
0726
0797
0623
06FA
05A1
04AB
0603
0209
0B48
1DDA
1E7E
1981
1830
14C1
130D
114A
0F85
0E60
0C64
0B43
09A1
07B1
0657
0511
0418
02FA
01DE
008D
FF74
FE82
FDAB
FCE1
FBD6
FB42
F97E
F8F4
F923
F764
F918
F320
E3AE
E110
E4B6
E480
E6C9
E773
E7FF
E9A1
E985
EA7F
EAF2
EBCA
ECF6
ED13
EE58
EEEB
EF70
F00D
F085
F217
F200
F25F
F385
F39E
F4B4
F4EB
F5A6
F6CF
F6BE
F7E3
F801
F81E
F911
F925
FA30
FA3E
FAA9
FB69
FB31
FC8F
FBF3
FCA4
FDD6
FC96
0019
F929
E827
E719
EC25
ED13
F022
F16E
F308
F51E
F621
F7FA
F8B5
FA3D
FBC5
FC65
FE21
FF06
000F
013B
01F4
0353
044D
04F8
05AF
06C6
0743
07EC
0958
0948
0A82
09DF
0B3B
17C8
1E23
1A84
1A7F
1930
17EA
17E4
1606
164A
1585
1489
1458
12CE
12CC
1248
1195
112B
1014
0FF6
0E94
0E40
0E87
0D01
0CDA
0C07
0B84
0B98
0A5F
09F8
0911
0907
08F9
07E2
0843
0713
06B0
06A1
0565
05DE
04D1
0507
046F
030D
04CA
00F7
0771
1AB2
1D31
17FA
167C
129F
1147
0F5E
0D43
0CB0
0A48
0909
0789
05E4
04B0
02F5
020C
0078
FF73
FE65
FCD1
FC66
FB60
FA85
F940
F86E
F802
F6A4
F728
F581
F59E
F4B6
E652
DDB8
E165
E180
E336
E551
E508
E6A3
E730
E803
E873
E8BF
EA3D
EA6F
EBA0
EC47
EC73
EE19
EE7C
EF3A
EFA0
EFD6
F11A
F169
F289
F329
F32E
F422
F46A
F5CA
F680
F680
F730
F6DC
F801
F869
F841
F985
F92E
FA4E
FA90
FA54
FC55
FAAF
FD13
FC5E
EBDC
E3E2
E93C
EB0C
ED5B
EFF9
F0ED
F314
F43C
F5A7
F74B
F845
F9BF
FAC2
FC03
FD89
FE57
FF8D
00F1
01BB
02E4
03D9
042D
056E
0623
06EA
07F5
0766
092E
0915
0961
1567
1D4C
1A38
19E3
187D
16D7
1770
15E4
1591
149E
13B7
1435
12B4
128A
1211
10DC
10EA
0FAC
0F43
0E9C
0D9A
0DC4
0CD7
0CC9
0C6A
0B5E
0B6F
0A7A
09D2
0918
089A
08A8
07A5
0781
06F9
06E0
06B1
0553
064E
0516
047A
056F
02D7
0466
02A0
02BE
150D
1F16
1943
1720
14CE
1232
10A9
0E27
0D3D
0B53
09C7
08D5
06DA
05B0
040D
02C4
020C
00C0
FF82
FE5A
FDA1
FC9A
FBE4
FAD6
F9AD
F94F
F7AA
F7AC
F6EF
F5B7
F737
ECF4
DF17
E020
E2C2
E33D
E5A4
E5D7
E712
E7F2
E81E
E97F
EA25
EB09
EB93
ECCD
EDB1
ED64
EECF
EF63
EFFF
F11D
F0E7
F1FC
F273
F2FB
F455
F462
F518
F552
F619
F749
F72F
F839
F848
F899
F978
F95B
FAFC
FAC0
FB02
FC39
FB8E
FD5C
FC4C
FD31
FE2E
EEFA
E4E7
EA1D
EBF2
EDEF
F0A1
F176
F41E
F549
F682
F7BE
F8AA
FAFC
FBF3
FCFC
FE65
FF67
00A7
0186
02AF
0390
04AD
057F
05F9
0755
078C
086D
095C
099F
09F0
08D2
110E
1D56
1CE8
1A7E
1A7E
1872
1860
176A
1698
1643
14FE
1504
13CB
1352
1339
11D6
120F
10F9
1027
1056
0EEA
0E8C
0DF8
0D70
0D44
0C80
0C7C
0B6C
0AAB
0A21
0951
09DA
08C8
0848
080C
0710
07B0
0648
05FA
0601
0492
05C4
03EE
043F
04DA
00F1
0DB0
1E01
1B9C
17C2
1603
12C1
11BA
0F56
0D82
0C5F
0AB7
0999
07A8
0603
0492
0385
02B2
011F
0065
FFD1
FE99
FD4F
FC41
FB4E
FA82
FA1A
F8D2
F896
F789
F641
F7DE
EEF0
E0DA
E0CA
E379
E387
E60A
E649
E70F
E80F
E832
E9C5
E9BD
EA14
EB6B
EC67
EDD5
ED92
EDB9
EEF7
EF5E
F023
F0C3
F1B4
F2F2
F382
F426
F490
F51F
F58B
F5F2
F6EE
F71D
F76F
F820
F876
F8EC
F939
FA33
FAD0
FA83
FB03
FB99
FC6A
FC9B
FC72
FD7A
FCC4
FBFB
FD39
FDE1
FE82
FF05
FF58
FFB4
FF9C
0016
0023
008B
0121
00EB
018F
019F
023A
02D5
024D
034F
0326
03B0
0475
0377
0500
037C
0490
061C
F84C
EE82
F05C
F586
039B
095A
0627
0806
06DF
06AA
07E4
069C
077C
06C4
06B4
07EA
0778
07FA
07C2
0859
08DB
07E8
082B
07E9
0813
0829
0774
07B4
076C
07DE
07E8
0772
082B
0790
0715
0730
073D
0774
06D6
0725
0732
06E4
071E
0669
0652
05D9
05CD
0690
05CC
05D6
05C3
054A
0584
04E4
04FD
04D9
04CF
0534
046F
04A7
049F
0454
0456
03B1
0414
0399
0363
03EF
0362
0396
029F
027D
0303
0241
032C
01E6
01C7
02F0
009B
0295
FF5F
F36C
EF85
F263
F49F
F371
F94A
0A09
0E38
09E8
0B00
0916
0826
084B
067A
06E7
05AD
04FB
057A
0406
0434
0418
033B
0328
025E
021A
0212
01B8
0144
00D5
00BF
FFFD
FF65
FF83
FF95
FF29
FE5F
FE5C
FE12
FDDF
FDFC
FD5B
FD9F
FD54
FC8F
FD10
FCA9
FC47
FC4D
FC1B
FC6E
FC41
FC13
FB7D
FB0C
FBA6
FBAC
FBE1
FBA0
FB2D
FB71
FAD3
FAF1
FADB
FA69
FAE5
FA65
FACF
FB26
FAAC
FAFD
FA50
FB04
FAB1
F9D5
FC36
F999
FBB6
0A79
0FAA
0B0C
0AC5
08D9
0674
06D0
04DE
042D
03E2
01D4
022A
FFC5
FF5C
00D7
F230
E3EC
E6BC
E8A8
E907
EB72
EB7B
ECE3
EDBD
EE6C
EFC7
EFCE
F0E2
F160
F1FB
F34C
F376
F44A
F49D
F4F8
F5F1
F64E
F713
F768
F810
F8FF
F96B
FA54
FA94
FB55
FBF5
FB95
FC1C
FC27
FCC6
FDE6
FDCC
FE55
FE91
FEA0
FF3A
FF66
001B
005A
0067
0121
0121
0160
0216
0241
0296
029F
0261
02EB
0334
031C
0349
038F
0460
03E5
04AD
0510
FB15
F26D
F52F
F6D9
F80B
FA55
FA2A
FBDE
FCC3
FD5A
FEE2
FF25
009F
00F6
01C4
034B
02AF
0409
04D2
0573
0651
060B
0881
069E
09DA
1A3E
1F3E
1AB1
1A8A
189D
175B
1697
14CE
1492
1370
12F1
1234
10A6
103B
0F05
0E71
0E02
0CC5
0C47
0B68
0AA9
0A4B
09F6
0970
0859
07ED
0732
064B
0598
043C
03F2
03D8
0349
02F4
0226
01C8
01BD
015F
00BB
005F
0063
FFA6
FFB7
FFC6
FECD
FEB8
FE5D
FDF4
FDC0
FD74
FDB5
FD10
FCDB
FD03
FC8B
FC8C
FBDF
FBEA
FC21
FBAA
FBFB
FBAD
FBAF
FB7E
FB47
FBCB
FABE
FB01
FB2F
FAB1
FB96
FB07
FB4D
FAD3
FA9A
FBE5
FA49
FB9C
FA22
FADC
09F2
104A
0CEC
0B61
0885
0973
FDA1
EBF4
ED72
EFFE
EFCD
F286
F195
F2B6
F376
F348
F4D1
F4D2
F582
F577
F5B3
F6D9
F6B1
F78A
F7C7
F813
F8EF
F903
F99C
F972
F9DD
FAB5
FAA1
FB5A
FBBC
FC41
FC8A
FC92
FD55
FD2B
FD6D
FDD6
FDE8
FEB2
FED1
FEFC
FF16
FF91
005D
FFDD
0003
005A
0080
00B4
0098
011B
00B6
0101
01BD
011F
01F0
01E2
01A8
0291
022A
0292
0299
0238
02A0
0282
0319
02CC
02D3
0349
02B4
0372
030F
032F
03AD
02E6
0410
031E
033F
0418
02CE
0591
FEB4
F298
F32B
F533
F731
F795
F9BA
0A1C
11FE
0D78
0DE0
0C89
0B98
0BF9
0A67
0AD9
0A06
0990
09C9
08A9
08BE
0810
07A5
0773
06D0
071A
0662
05ED
05A9
0559
0598
0498
045B
0442
03C1
03EE
0308
02BB
0297
0232
0288
0220
0203
01C2
015F
0172
00EE
0104
009F
004C
0087
0008
003B
FFFA
FFB5
FFD2
FF66
FFC1
FF4A
FF41
FF8A
FE9D
FEF7
FEB7
FE72
FEAD
FE20
FE88
FE2C
FE21
FE7D
FDF4
FE5D
FDD0
FDDF
FDFD
FD80
FE1C
FD58
FE2D
FE2C
FD0C
FE5D
FD1A
FE59
FD88
FD0E
0B4C
12D2
0F60
0E3E
0B99
0C75
024C
EFF2
EFE8
F2C5
F201
F4C6
F491
F56F
F607
F5BA
F70F
F6C2
F780
F7D0
F7BB
F8C2
F8BA
F99D
F9ED
F9D8
FAA2
FADA
FB76
FB7B
FBA0
FC25
FC2A
FCD8
FCD4
FD26
FDB8
FDC6
FE3A
FDD2
FE38
FEF1
FECA
FF52
FF37
FF89
000D
FFD4
001D
FFF2
003D
0084
0069
00DC
00A7
00FE
012D
00FF
019C
0157
0194
01D3
01B6
022C
01D1
0201
0215
01DE
0242
01EE
0234
0214
01E9
0239
01D5
0299
0245
022B
02E2
021F
02D7
01FF
0208
0303
011E
03CD
FEB8
F20D
F1A8
F3E4
F54D
F62A
F74E
06AE
1080
0C23
0C40
0B5E
09A2
0A3A
08DD
08D1
0834
07D4
07FE
06D5
0700
065A
05DC
05CF
0505
0546
048A
03F1
03DA
0321
0325
02A9
029F
0293
0203
0240
0195
011F
0115
00D4
00BB
000C
001F
FFF8
FF8A
FFCA
FF58
FF5C
FF25
FEE3
FF01
FE73
FE89
FE2D
FE12
FE4F
FD84
FDF0
FDC8
FD68
FDD9
FD57
FD7E
FD21
FD0D
FD74
FCBC
FD22
FCE9
FCD9
FD4F
FC7D
FD1A
FCFF
FCBE
FCFE
FC6D
FD20
FC7B
FC98
FCF0
FBE6
FD43
FC32
FCDB
FD00
FB28
082B
1231
0E98
0DF4
0ABD
0AD1
0739
F3D8
ED03
F189
F0E8
F2CC
F3ED
F407
F548
F521
F5E1
F616
F6A1
F742
F6FA
F7DA
F83B
F8C5
F922
F929
FA27
FA40
FAC1
FB23
FADE
FBC1
FBDB
FC16
FCA5
FCAC
FD51
FD74
FD9C
FDEE
FE1D
FED3
FEF2
FF09
FF2C
FF3F
FFA8
FFAA
FFF6
0026
004B
00B7
00D1
0123
0103
0129
01AA
017E
01E1
01E7
01F8
024B
01EC
0230
0220
024E
02EA
027A
028B
02B5
0302
0324
02C2
0312
02C9
031E
034F
02D9
0342
02D5
038C
0378
02FD
0424
028E
045B
00EB
F3B0
F1FB
F4C7
F58E
F85F
F6E7
019D
1095
0EE6
0D5F
0DAB
0B33
0B84
0A82
0A1C
0A04
0901
0950
0889
0825
07E7
076A
075E
06A2
066B
05D1
0572
0581
04D6
04E3
044A
03E4
0402
035E
0378
0301
0288
0286
0215
0226
01B6
018D
019F
0133
0159
00FC
00E3
00AB
0034
0082
FFFC
FFC8
FFB7
FF5C
FF8F
FF0C
FF41
FF34
FE9B
FF06
FEA4
FE87
FE50
FDE7
FE6E
FE03
FDF2
FE24
FE12
FE2F
FDA4
FDFD
FDDA
FDC7
FE19
FD7F
FE31
FDCA
FD88
FDDF
FCED
FE25
FD58
FDD3
FE59
FBAA
0774
1308
0FA0
0EC3
0BED
0B52
0980
F670
EDA7
F288
F19E
F34B
F4DE
F46F
F5DD
F5C5
F68A
F6E1
F725
F80B
F7DC
F8CF
F903
F927
F9C8
F9BE
FAD1
FB07
FB22
FBD9
FBD4
FC5F
FC72
FCB7
FCF1
FCFD
FE0D
FE32
FE88
FEE8
FEA6
FF25
FF38
FFBA
FFE4
FFAB
0063
0045
00A6
00E4
00A3
0122
00FB
0138
0151
018E
021C
0183
0236
024C
01E5
0292
0240
02DD
02EF
0299
030C
024C
02EA
0313
02C9
0362
02BA
0379
036D
02EC
0369
02B1
0352
0300
02D0
033E
02A7
03F3
0242
039E
0244
F469
F139
F4B1
F450
F7C7
F68B
FE88
0D40
0CBF
0BA8
0B96
0938
09AB
086B
0925
07DC
07B9
0841
FB12
F2B5
F66E
F717
F8B9
FA1D
F9F5
FB68
FBAF
FCA3
FD66
FDB9
FEE6
FF34
FFA9
002B
00B0
013B
018B
026A
02AC
02CB
033D
0390
0450
0440
0404
0472
04AE
0521
05A8
05B2
05AA
05E8
05E9
05FA
0664
0635
0626
0634
0628
06A0
0649
0609
067F
063B
0625
0673
063F
05CD
0607
0636
057F
05AF
05B5
050F
0554
054F
0538
04DB
049F
04F7
0448
04AC
0464
03CF
04B8
0232
06CB
1391
150F
113E
10D3
0E60
0D1D
0C0F
0A43
09E3
0871
0789
06FA
0585
04D7
040B
031E
0217
011E
00AE
FFF4
FF4B
FE68
FD6C
FCE4
FC74
FC19
FB5E
FAB8
FA45
F9BD
F952
F8AE
F8B3
F864
F786
F7BC
F733
F647
F664
F65A
F60A
F584
F57C
F595
F513
F50C
F50F
F4D7
F47D
F416
F420
F40E
F438
F475
F445
F40C
F3DE
F43C
F459
F434
F438
F3F0
F44A
F488
F46F
F4AE
F4C3
F521
F4F8
F507
F595
F559
F5C4
F5E9
F5B4
F5D2
F5AF
F663
F623
F64A
F717
F665
F770
F73C
F7C8
F8C3
EE71
E5AB
E8C4
EAB8
EC18
EE5B
EEF5
F0C1
F19E
F287
F3FC
F480
F614
F70A
F782
F8C7
F99C
FAA1
FB6E
FBF4
FCA7
FD60
FE71
FF29
FFA9
0039
00B0
016D
0223
02D2
0326
036B
0453
04ED
0543
05A0
05C0
063A
06C8
06EC
0743
07DB
07EF
0811
08A9
089F
08B2
0944
094B
094E
098D
09C3
09E1
09ED
0A1D
0A00
0A0D
0A65
0A41
0A36
0A8E
0AAB
0A55
0A23
0A12
09ED
0A46
0A43
0A26
0A73
0A24
0A33
0A15
09A1
09D0
097E
09C3
09C5
0901
0961
0918
08E1
0878
0843
094B
06E9
0A92
1708
19DD
15FD
14FE
12EA
11AD
10E7
0F4F
0EC0
0DC8
0CAA
0B5D
0A4D
09F0
08D9
07FD
0741
066D
05D9
04DE
0431
03C6
032C
0228
0153
014B
00A8
FFEB
FF5F
FE89
FE48
FDF1
FDA1
FD43
FC7A
FC41
FC08
FBA0
FB5A
FB5B
FB7D
FAE3
FA60
FA1B
F9ED
F9E6
F9AD
F9DF
F979
F932
F9CE
F94A
F8D1
F8E7
F8D8
F911
F8EC
F8B5
F863
F8B3
F936
F8B9
F90D
F919
F8B5
F8FF
F8B4
F913
F910
F8BC
F953
F92B
F97E
F977
F94C
F9FC
F9A9
FA1B
FA04
F9F2
FAE1
FA17
FB10
FAA3
FA70
FC9C
F34C
E93B
EB65
ED56
EECA
F0CA
F1B7
F35E
F3CA
F5B4
F50D
F7E5
05C6
0AFF
07C4
089B
0780
069D
06DE
062B
06A0
05C8
0593
05FF
0567
05C8
0555
04DC
04F0
0490
04A1
0413
03ED
0442
0400
0415
03DC
03C0
03B9
0349
0336
02FD
032B
0352
02E6
02CD
0291
0272
0268
024A
0267
024F
0243
01E2
01E0
027E
0236
0213
0216
01CD
01FA
01EB
01DC
01CF
0191
017C
0149
0188
019A
016A
0186
0160
017B
015E
0142
01B6
016E
012C
0125
00F3
013A
0150
0151
0134
011A
015E
0116
00D6
00FB
012E
0156
0106
0102
0113
0108
012E
00F4
0109
0131
00F8
00EE
00CE
0103
011C
00C1
00BC
00AD
00DD
010F
00F9
00FD
00A4
00B9
00F9
00A3
00D5
00CB
007F
00DB
00DD
00A3
0091
0079
00C2
00F4
00BF
00A9
00C5
00AC
006F
0064
0066
006C
0073
0074
00A5
00B1
0083
0073
0051
0052
006A
001D
0021
006B
0030
001F
003A
000D
000E
0025
0047
0046
0011
0037
001E
FFD6
FFFC
FFFB
0016
0033
FFF5
FFF3
FFDE
FFBD
FFE8
FFD1
FFB3
FFE3
FFEF
FF99
FF87
FFDA
FF94
FF4A
FF8A
FF71
FF78
FFAD
FF7F
FF78
FF60
FF3F
FF66
FF4C
FF43
FF4E
FF32
FF45
FF34
FF33
FF48
FF0E
FF13
FF05
FEC6
FEF8
FF03
FEFC
FF23
FEEB
FED0
FEEF
FECF
FEB6
FEBC
FEAC
FE9C
FEBC
FEBD
FE81
FE88
FE9D
FE7D
FE86
FEAB
FEA6
FE92
FE9B
FE91
FE76
FE88
FE83
FE64
FE60
FE5B
FE74
FE89
FE65
FE4C
FE4F
FE4C
FE4F
FE69
FE6F
FE49
FE3B
FE53
FE4B
FE27
FE34
FE57
FE4E
FE3F
FE3F
FE40
FE34
FE28
FE50
FE46
FE1B
FE3E
FE21
FE0A
FE3D
FE21
FE14
FE1B
FE1D
FE40
FE16
FE1D
FE57
FE43
FE71
FE85
FE45
FE45
FE44
FE50
FE70
FE50
FE4E
FE62
FE4F
FE52
FE5E
FE63
FE76
FE6F
FE68
FE8A
FE7D
FE66
FE82
FE8A
FEA0
FE9D
FE62
FE74
FE7D
FE6D
FE9E
FEA0
FE97
FEB3
FEBD
FECF
FEBD
FEC0
FEEB
FEDA
FEE2
FEFB
FED8
FEDA
FEFA
FEFB
FEF6
FF00
FF11
FF05
FEF9
FF19
FF2F
FF1E
FF29
FF4A
FF3C
FF29
FF35
FF41
FF50
FF5E
FF67
FF67
FF5F
FF6F
FF7C
FF83
FF92
FF90
FF94
FFA0
FF9F
FFA8
FFAA
FFA7
FFAE
FFBA
FFC2
FFC5
FFD9
FFE7
FFDD
FFE6
FFFA
FFFF
0001
0009
0013
0018
0025
002C
002A
0031
002F
0038
004C
004F
0058
005D
005E
0069
006A
0074
0080
007F
008A
008B
008E
00A0
00A4
00A7
00A8
00AB
00BA
00BA
00BC
00CE
00D4
00D3
00D8
00E2
00E6
00EA
00F8
00F8
00F6
0100
0103
010A
0111
0112
0119
011D
0123
012B
012B
0133
0137
0138
013F
0142
0148
014E
014F
0154
0155
0158
0160
0161
0164
0169
016F
016F
0171
017A
0177
017A
017F
0180
018A
0186
0186
018D
018B
0192
018D
0193
0199
0190
019D
019A
019C
01A1
0197
01AC
019A
01A4
01AF
017D
0235
0312
02D8
02B4
02B1
027C
027F
0268
0253
024D
0234
022D
021A
0210
0201
01EA
01EB
01D4
01C9
01C4
01AE
01AB
019C
0191
018B
017B
0179
016C
0162
015A
014D
014C
013D
0138
0137
0128
0124
011A
0114
0110
0106
0108
00FD
00F6
00F5
00EB
00EB
00E4
00DF
00DD
00D4
00D6
00D0
00C9
00C9
00C4
00C3
00BD
00B9
00B9
00B5
00B4
00AE
00AC
00AD
00A8
00A7
00A3
00A1
00A1
009A
009B
009C
0098
0093
0092
0093
008E
008E
008D
0087
008A
0089
0085
0085
0084
0080
007D
007E
007D
007B
0079
0076
0078
0075
0072
0074
0070
006C
006E
006C
0067
0066
0066
0061
0061
0060
005C
005D
005A
0058
0057
0051
004F
0050
004E
004D
004A
0047
0044
0041
003F
003E
003C
0038
0036
0034
0031
002E
002A
002A
0026
0022
0022
001C
001B
001A
0015
0014
0010
000B
0009
0006
0006
0001
FFFC
FFFC
FFF6
FFF3
FFF0
FFED
FFED
FFE7
FFE3
FFE2
FFDC
FFD9
FFD7
FFD1
FFD1
FFCD
FFC6
FFC6
FFC3
FFBE
FFBA
FFB6
FFB6
FFB4
FFAB
FFA8
FFA6
FFA2
FFA0
FF9D
FF98
FF95
FF91
FF8F
FF8B
FF86
FF85
FF83
FF7D
FF78
FF74
FF71
FF70
FF6E
FF66
FF64
FF64
FF5F
FF5B
FF59
FF56
FF52
FF4F
FF4D
FF49
FF47
FF44
FF3F
FF3F
FF3C
FF36
FF35
FF32
FF30
FF2A
FF27
FF2B
FF25
FF1F
FF20
FF1D
FF1A
FF17
FF13
FF13
FF11
FF0F
FF0C
FF08
FF08
FF04
FF03
FF03
FEFF
FEFE
FEFD
FEF9
FEF7
FEF8
FEF5
FEF2
FEF3
FEF0
FEED
FEF0
FEED
FEEA
FEEA
FEE7
FEE8
FEE7
FEE5
FEE5
FEE2
FEE1
FEE4
FEDF
FEDE
FEE1
FEDE
FEDC
FEDF
FEDD
FEDC
FEDD
FEDB
FEDC
FEDC
FEDB
FEDD
FEDA
FEDA
FEDD
FEDB
FEDB
FEDD
FEDC
FEDC
FEDF
FEDF
FEDE
FEE0
FEE0
FEDF
FEE2
FEE3
FEE4
FEE5
FEE6
FEE6
FEE7
FEE9
FEEB
FEEC
FEEE
FEEE
FEEF
FEF3
FEF2
FEF2
FEF7
FEF9
FEF9
FEFB
FEFD
FEFF
FF00
FF03
FF05
FF06
FF09
FF0B
FF0D
FF0F
FF12
FF14
FF16
FF19
FF1B
FF1D
FF20
FF23
FF24
FF27
FF2A
FF2D
FF30
FF32
FF34
FF37
FF3B
FF3D
FF40
FF43
FF46
FF4A
FF4C
FF4F
FF52
FF55
FF58
FF5C
FF5E
FF61
FF65
FF68
FF6B
FF6E
FF72
FF75
FF78
FF7C
FF7F
FF82
FF86
FF8A
FF8C
FF90
FF93
FF96
FF9A
FF9D
FFA1
FFA4
FFA7
FFAB
FFAE
FFB2
FFB5
FFB8
FFBC
FFBF
FFC3
FFC6
FFCA
FFCD
FFD1
FFD5
FFD8
FFDC
FFDF
FFE2
FFE6
FFE9
FFED
FFF1
FFF4
FFF7
FFFB
FFFE
0001
0005
0008
000B
000F
0012
0016
0019
001C
001F
0023
0026
0029
002C
0030
0033
0036
003A
003D
003F
0043
0046
0048
004C
004F
0052
0055
0057
005B
005D
0060
0063
0066
0069
006C
006E
0071
0074
0076
0079
007B
007E
0080
0083
0085
0088
008A
008D
008F
0091
0094
0095
0098
009A
009B
009E
00A1
00A2
00A4
00A6
00A8
00AA
00AB
00AE
00AF
00B1
00B3
00B4
00B6
00B8
00B8
00BB
00BC
00BD
00BF
00C0
00C1
00C2
00C4
00C5
00C6
00C8
00C8
00C9
00CB
00CB
00CC
00CE
00CE
00CF
00CF
00D0
00D1
00D1
00D2
00D2
00D3
00D5
00D4
00D4
00D5
00D4
00D6
00D6
00D6
00D6
00D6
00D6
00D7
00D7
00D6
00D6
00D6
00D6
00D6
00D6
00D5
00D6
00D5
00D5
00D4
00D3
00D4
00D3
00D3
00D2
00D1
00D1
00D0
00CF
00CF
00CD
00CD
00CC
00CA
00CB
00CA
00C8
00C8
00C7
00C6
00C4
00C3
00C3
00C1
00C0
00BF
00BE
00BC
00BB
00BA
00B8
00B7
00B5
00B4
00B3
00B0
00AF
00AF
00AB
00AB
00AA
00A6
00A6
00A5
00A2
00A1
009E
009D
009B
0099
0098
0096
0094
0092
0090
008F
008C
008A
0089
0086
0084
0083
0081
007E
007D
007B
0078
0077
0075
0071
0071
006E
006B
006B
0067
0065
0064
0060
005F
005D
005A
0058
0055
0053
0052
004F
004D
004B
0048
0046
0044
0041
003F
003D
003B
0039
0035
0035
0032
002E
002D
002B
0029
0027
0023
0022
0021
001D
001B
0019
0017
0014
0013
0011
000E
000C
000A
0008
0006
0002
0001
FFFF
FFFC
FFFB
FFF9
FFF6
FFF4
FFF3
FFF1
FFED
FFEC
FFEA
FFE8
FFE6
FFE3
FFE3
FFE1
FFDE
FFDD
FFDA
FFD8
FFD7
FFD5
FFD3
FFD2
FFCF
FFCD
FFCC
FFCB
FFC8
FFC6
FFC5
FFC3
FFC1
FFC0
FFBE
FFBD
FFBB
FFB9
FFB8
FFB6
FFB5
FFB4
FFB1
FFB0
FFAF
FFAE
FFAC
FFAA
FFA9
FFA9
FFA6
FFA4
FFA4
FFA2
FFA1
FFA0
FF9F
FF9E
FF9D
FF9B
FF9A
FF99
FF98
FF97
FF96
FF95
FF94
FF94
FF92
FF91
FF91
FF8F
FF8F
FF8E
FF8D
FF8C
FF8C
FF8B
FF8A
FF8A
FF89
FF88
FF88
FF87
FF86
FF87
FF85
FF84
FF84
FF84
FF84
FF83
FF81
FF82
FF83
FF81
FF81
FF82
FF80
FF80
FF81
FF80
FF80
FF80
FF80
FF80
FF7F
FF7F
FF80
FF7F
FF7F
FF80
FF7F
FF80
FF80
FF80
FF80
FF80
FF80
FF81
FF81
FF82
FF81
FF81
FF83
FF82
FF82
FF84
FF83
FF84
FF86
FF85
FF85
FF87
FF87
FF86
FF88
FF88
FF88
FF8A
FF8A
FF8A
FF8B
FF8C
FF8C
FF8D
FF8E
FF8E
FF8F
FF90
FF91
FF92
FF92
FF93
FF94
FF95
FF96
FF97
FF98
FF98
FF9A
FF9B
FF9A
FF9C
FF9E
FF9E
FFA0
FFA0
FFA1
FFA3
FFA3
FFA4
FFA6
FFA6
FFA8
FFA9
FFA9
FFAC
FFAB
FFAD
FFAF
FFAF
FFB0
FFB1
FFB3
FFB5
FFB4
FFB6
FFB8
FFB8
FFBA
FFBB
FFBC
FFBD
FFC0
FFC0
FFC1
FFC3
FFC4
FFC5
FFC7
FFC7
FFC9
FFCB
FFCC
FFCD
FFCD
FFCF
FFD1
FFD2
FFD3
FFD4
FFD6
FFD7
FFD8
FFDB
FFDB
FFDC
FFDF
FFDF
FFE0
FFE2
FFE3
FFE4
FFE6
FFE7
FFE8
FFEA
FFEA
FFEC
FFED
FFED
FFF0
FFF1
FFF2
FFF3
FFF4
FFF6
FFF6
FFF9
FFF9
FFFA
FFFC
FFFD
FFFE
FFFF
0000
0002
0002
0005
0006
0005
0008
0009
000A
000B
000B
000E
000E
000F
0011
0011
0013
0013
0015
0017
0016
0019
0019
001A
001C
001B
001E
001F
001F
0020
0021
0022
0023
0024
0025
0025
0027
0027
0028
002A
002A
002B
002C
002D
002E
002E
0030
0030
0030
0031
0031
0034
0033
0033
0036
0035
0036
0038
0037
0038
0039
0039
003A
003A
003B
003C
003C
003C
003D
003D
003D
003F
003E
003F
0040
003F
0040
0041
0041
0042
0041
0043
0043
0042
0044
0043
0043
0045
0044
0045
0045
0045
0046
0045
0046
0046
0045
0046
0047
0046
0046
0047
0046
0047
0047
0047
0047
0046
0047
0048
0046
0047
0047
0046
0047
0047
0046
0047
0045
0045
0046
0045
0045
0045
0045
0045
0045
0044
0044
0044
0044
0044
0043
0043
0043
0041
0042
0043
0041
0040
0041
0040
0040
003F
003F
003F
003F
003E
003D
003D
003D
003B
003C
003C
003B
003A
003A
003A
0039
0039
0038
0037
0037
0036
0036
0036
0034
0035
0034
0033
0033
0032
0032
0031
0030
0030
002F
002F
002E
002D
002D
002C
002B
002B
002A
002A
0029
0028
0028
0027
0026
0025
0025
0025
0023
0023
0023
0021
0021
0021
001F
001E
001F
001D
001C
001D
001B
001B
001B
0018
0019
0018
0016
0017
0016
0014
0014
0014
0013
0013
0011
0011
0011
000F
000F
000E
000E
000D
000C
000B
000B
000A
0009
0008
0008
0007
0006
0006
0005
0005
0004
0003
0003
0002
0001
0000
0000
0000
FFFE
FFFE
FFFE
FFFC
FFFC
FFFC
FFFA
FFFA
FFFA
FFF9
FFF8
FFF8
FFF7
FFF7
FFF7
FFF5
FFF5
FFF5
FFF3
FFF3
FFF3
FFF2
FFF2
FFF1
FFF0
FFF0
FFEF
FFEF
FFEF
FFED
FFEE
FFED
FFEC
FFEC
FFEB
FFEB
FFEB
FFE9
FFEA
FFEA
FFE8
FFE8
FFE9
FFE7
FFE6
FFE7
FFE7
FFE6
FFE6
FFE5
FFE6
FFE4
FFE3
FFE4
FFE4
FFE3
FFE3
FFE2
FFE2
FFE2
FFE1
FFE2
FFE0
FFE0
FFE1
FFDF
FFDF
FFE0
FFDE
FFDF
FFDF
FFDE
FFDE
FFDD
FFDE
FFDE
FFDC
FFDE
FFDD
FFDC
FFDD
FFDD
FFDC
FFDC
FFDC
FFDC
FFDB
FFDC
FFDB
FFDB
FFDC
FFDC
FFDB
FFDB
FFDC
FFDB
FFDA
FFDB
FFDB
FFDA
FFDA
FFDA
FFDB
FFDA
FFD9
FFDC
FFDA
FFDA
FFDB
FFDA
FFDB
FFDB
FFDA
FFDB
FFDB
FFDB
FFDB
FFDB
FFDB
FFDB
FFDB
FFDB
FFDC
FFDC
FFDC
FFDC
FFDB
FFDD
FFDC
FFDC
FFDD
FFDC
FFDD
FFDD
FFDD
FFDD
FFDD
FFDE
FFDE
FFDD
FFDF
FFDF
FFDE
FFDF
FFDF
FFDF
FFDF
FFDF
FFE0
FFE0
FFE0
FFE0
FFE0
FFE1
FFE1
FFE1
FFE1
FFE3
FFE2
FFE1
FFE3
FFE4
FFE3
FFE4
FFE5
FFE4
FFE5
FFE5
FFE4
FFE6
FFE6
FFE5
FFE7
FFE7
FFE6
FFE7
FFE8
FFE8
FFE7
FFE9
FFEA
FFE8
FFEA
FFEA
FFEA
FFEB
FFEA
FFEB
FFEC
FFEC
FFED
FFEB
FFEE
FFEF
FFED
FFEE
FFEF
FFEF
FFF0
FFEF
FFF0
FFF0
FFF0
FFF1
FFF2
FFF2
FFF2
FFF3
FFF2
FFF4
FFF4
FFF3
FFF5
FFF5
FFF5
FFF6
FFF5
FFF7
FFF7
FFF7
FFF8
FFF8
FFF8
FFF9
FFF8
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFD
FFFC
FFFC
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0001
0002
0000
0002
0003
0002
0004
0004
0003
0005
0004
0005
0006
0005
0006
0006
0006
0007
0007
0007
0008
0008
0008
0008
000A
0009
0008
000A
000A
0009
000B
000A
000A
000B
000B
000D
000B
000B
000E
000C
000C
000E
000D
000D
000E
000D
000E
000E
000E
000F
000F
000E
000F
0010
000F
000F
0010
000F
0011
0010
0010
0011
0010
0011
0011
0011
0011
0011
0012
0011
0011
0013
0011
0012
0013
0012
0012
0013
0013
0012
0012
0014
0013
0013
0013
0013
0013
0013
0014
0014
0013
0014
0014
0013
0014
0014
0014
0014
0014
0013
0014
0014
0014
0014
0014
0014
0014
0013
0015
0015
0013
0014
0014
0014
0014
0013
0014
0014
0013
0014
0013
0014
0014
0013
0014
0013
0012
0014
0013
0013
0013
0013
0013
0012
0013
0012
0012
0012
0012
0013
0012
0012
0012
0010
0012
0012
0010
0011
0011
0011
0011
0010
0011
0010
0010
0011
0010
0010
000F
0010
0010
000F
0010
000F
000E
0010
000E
000E
000F
000E
000E
000E
000D
000D
000D
000C
000D
000C
000C
000C
000C
000B
000C
000C
000B
000B
000B
000B
000A
000B
000A
000A
000B
0009
0009
000A
0008
000A
0008
0008
0009
0007
0008
0008
0007
0007
0006
0007
0007
0006
0007
0007
0005
0006
0006
0005
0005
0006
0004
0005
0004
0003
0005
0004
0002
0004
0003
0003
0003
0002
0003
0002
0001
0002
0002
0001
0001
0001
0001
0000
0001
FFFF
0000
0000
FFFF
0000
FFFE
FFFE
0000
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFA
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFA
FFF8
FFF9
FFF9
FFF8
FFFA
FFF8
FFF8
FFF9
FFF7
FFF8
FFF8
FFF7
FFF9
FFF7
FFF8
FFF8
FFF6
FFF8
FFF7
FFF7
FFF8
FFF7
FFF7
FFF7
FFF7
FFF7
FFF7
FFF7
FFF6
FFF7
FFF7
FFF5
FFF8
FFF7
FFF5
FFF7
FFF6
FFF6
FFF6
FFF5
FFF6
FFF6
FFF5
FFF6
FFF6
FFF6
FFF5
FFF6
FFF6
FFF5
FFF6
FFF5
FFF5
FFF7
FFF5
FFF5
FFF6
FFF5
FFF6
FFF6
FFF4
FFF5
FFF6
FFF5
FFF5
FFF5
FFF5
FFF6
FFF6
FFF5
FFF6
FFF6
FFF5
FFF6
FFF6
FFF5
FFF7
FFF6
FFF5
FFF6
FFF6
FFF6
FFF6
FFF6
FFF6
FFF5
FFF5
FFF6
FFF5
FFF6
FFF7
FFF6
FFF5
FFF7
FFF6
FFF6
FFF7
FFF6
FFF7
FFF6
FFF7
FFF8
FFF6
FFF7
FFF8
FFF6
FFF7
FFF7
FFF7
FFF7
FFF7
FFF8
FFF7
FFF8
FFF8
FFF7
FFF9
FFF8
FFF7
FFF9
FFF7
FFF8
FFF9
FFF8
FFF9
FFF9
FFF9
FFF8
FFF8
FFFA
FFF8
FFF9
FFF9
FFF8
FFFA
FFF8
FFF9
FFFB
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFC
FFFB
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFD
FFFC
FFFC
FFFD
FFFC
FFFD
FFFE
FFFD
FFFE
FFFE
FFFD
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0001
0001
0001
0001
0002
0001
0001
0002
0002
0001
0001
0002
0002
0001
0002
0002
0002
0002
0002
0003
0003
0003
0002
0003
0004
0002
0003
0004
0003
0002
0004
0003
0002
0005
0004
0003
0004
0003
0004
0004
0003
0005
0004
0004
0005
0004
0005
0005
0004
0005
0004
0005
0005
0003
0005
0005
0005
0005
0005
0005
0005
0006
0005
0005
0005
0005
0006
0005
0004
0006
0005
0005
0006
0004
0005
0006
0005
0005
0005
0005
0005
0005
0005
0005
0006
0005
0005
0006
0006
0005
0005
0007
0005
0005
0007
0005
0005
0006
0005
0005
0006
0005
0006
0006
0006
0005
0006
0006
0005
0006
0006
0006
0006
0006
0005
0006
0006
0006
0005
0006
0005
0005
0006
0005
0005
0005
0005
0006
0005
0005
0006
0005
0005
0005
0005
0006
0004
0006
0005
0003
0007
0005
0003
0005
0005
0005
0005
0005
0006
0004
0005
0006
0004
0005
0005
0004
0005
0004
0004
0005
0004
0004
0004
0004
0005
0004
0004
0004
0004
0004
0003
0003
0004
0004
0003
0004
0004
0003
0004
0003
0003
0003
0003
0003
0003
0003
0002
0002
0003
0003
0003
0002
0002
0003
0002
0002
0002
0002
0003
0002
0002
0002
0001
0003
0002
0001
0002
0002
0002
0002
0001
0002
0001
0001
0002
0001
0001
0001
0001
0000
0001
0001
0000
0001
0001
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFE
0000
0000
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFD
FFFF
FFFD
FFFE
FFFF
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFE
FFFD
FFFE
FFFE
FFFD
FFFE
FFFD
FFFD
FFFF
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFC
FFFE
FFFD
FFFD
FFFE
FFFC
FFFD
FFFD
FFFD
FFFE
FFFC
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFE
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFC
FFFE
FFFF
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
FFFE
FFFF
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
0001
FFFF
0000
0001
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0001
0000
0000
0001
0001
0000
0000
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0002
0001
0000
0001
0002
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0002
0000
0001
0002
0000
0002
0001
0001
0002
0000
0002
0001
0001
0002
0000
0002
0002
0000
0002
0002
0001
0002
0002
0002
0001
0002
0002
0001
0002
0001
0002
0002
0001
0002
0001
0001
0002
0001
0001
0002
0001
0001
0002
0001
0002
0001
0001
0002
0001
0001
0002
0002
0001
0002
0002
0002
0001
0002
0002
0002
0002
0002
0002
0002
0001
0002
0002
0002
0002
0001
0002
0003
0001
0002
0002
0001
0002
0001
0002
0002
0001
0003
0001
0001
0002
0000
0002
0002
0001
0002
0001
0002
0002
0000
0002
0002
0001
0002
0001
0001
0001
0001
0002
0001
0002
0001
0000
0003
0001
0001
0002
0000
0002
0002
0000
0002
0001
0000
0001
0001
0001
0001
0000
0001
0002
0000
0001
0001
0001
0001
0000
0002
0001
0000
0002
0001
0000
0002
0000
0001
0002
0000
0001
0000
0001
0001
0000
0001
0001
0000
0001
0000
0001
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
FFFF
0001
0001
FFFF
0001
0001
0000
0001
FFFF
0001
0001
0000
0000
FFFF
0001
0001
FFFF
0002
0000
FFFF
0001
FFFF
0000
0000
FFFF
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0001
FFFF
FFFF
0001
FFFF
0000
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFE
FFFF
0000
FFFE
FFFF
0000
FFFF
FFFE
0000
FFFF
FFFF
0000
FFFF
FFFE
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
0000
0000
FFFF
FFFF
0000
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
0001
FFFF
FFFF
0000
FFFF
FFFF
0001
FFFF
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0002
0000
0000
0002
0000
0000
0001
0000
0001
0000
0001
0001
FFFF
0001
0000
0000
0002
0000
0000
0001
0000
0000
0000
0001
0001
FFFF
0001
0001
FFFF
0001
0001
0001
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0001
0000
0000
0001
0001
0000
0001
0002
0000
0000
0002
0000
0000
0001
0001
0001
0001
0000
0001
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0001
0000
0000
0001
0000
0000
0001
0000
0001
0001
FFFF
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0001
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0001
0001
0000
0001
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0001
0000
0000
0002
0000
0000
0001
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0001
0001
FFFE
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
0001
0000
0000
0001
0000
FFFF
0001
0001
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFE
0000
0001
FFFF
0000
0001
0000
0000
0001
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0001
0000
0000
0001
FFFF
0000
0001
0000
0001
0000
0000
0001
0000
0000
0001
0000
0001
0000
0000
0001
0000
0000
0001
FFFF
0001
0001
0000
0001
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0001
0000
0000
0002
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0001
0000
FFFF
0001
0001
FFFF
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
FFFF
0001
0000
0000
0001
FFFF
0000
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFE
0001
0000
FFFE
0002
0001
FFFF
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0000
0000
0000
FFFF
0001
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0001
FFFF
0000
0000
0000
0001
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
FFFF
0000
0001
0000
0001
0000
FFFF
0001
0000
FFFF
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
FFFF
0000
0001
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
FFFF
0001
0000
FFFF
0001
0000
FFFF
0001
0001
FFFF
0001
0001
0000
0001
0001
0000
0001
0000
0000
0001
0000
0001
0000
0000
0001
0000
0001
0000
FFFF
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
FFFF
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0000
0001
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
FFFF
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0001
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0001
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0001
FFFF
FFFF
0000
0000
0000
0000
0001
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0001
0000
0000
0001
0000
0001
0000
0000
0000
0001
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0001
0000
FFFF
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
FFFF
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0002
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
FFFF
0001
0001
FFFE
0001
0000
FFFE
0001
0000
0000
0000
FFFF
0001
FFFF
0000
0001
FFFF
0001
0001
0000
0000
0001
0000
0000
0001
0000
FFFF
0002
FFFF
0000
0001
FFFF
0001
0000
0000
0001
FFFF
0001
0000
FFFF
0001
0000
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0001
0000
0001
0001
FFFF
0000
0001
FFFF
FFFF
0001
0000
FFFF
0000
FFFF
0000
0001
FFFE
0000
0001
FFFF
0001
0001
FFFF
0001
0000
0000
0001
0000
0001
0001
FFFF
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0000
0000
0000
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0001
0000
FFFF
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
FFFF
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
FFFF
0000
0000
FFFF
0001
0000
0000
0001
FFFF
0001
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
FFFF
FFFF
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0001
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0001
FFFF
0000
0000
FFFF
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0001
FFFF
0000
0000
0000
0001
0001
0000
0001
0000
0000
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0001
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0001
FFFF
0000
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
FFFF
0000
0001
0000
0000
0000
0000
0001
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0000
FFFF
0000
0001
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
FFFF
0000
0000
FFFF
0001
0001
FFFF
0000
0001
0001
0000
0000
0001
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0001
0001
FFFE
0000
0001
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0000
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0002
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0001
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0001
FFFF
0000
0001
0001
0000
0000
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0001
FFFF
FFFF
0001
0000
0000
FFFF
0000
0001
FFFF
0000
0000
FFFE
0000
0001
FFFF
0000
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0001
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
FFFF
0001
0000
FFFE
0000
0001
FFFF
0001
0000
FFFF
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
0000
0000
FFFF
0000
0000
FFFF
0001
FFFF
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0001
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0001
0000
FFFF
0001
0001
FFFF
0001
0001
FFFF
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0001
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0000
FFFF
0000
0000
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0001
0000
0001
0001
0001
0001
0000
0001
0002
0000
0001
0002
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
FFFF
0000
0002
0000
0001
0001
0000
0001
0000
0000
0001
0000
0001
0001
0000
0001
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0001
0001
0000
0001
0001
0001
0000
0000
0001
0000
0000
0001
0001
0001
0001
0001
0000
0002
0001
0000
0001
0000
0001
0002
0001
0001
0001
0001
0001
0000
0001
0000
0000
0002
0000
0000
0001
0000
0001
0001
0000
0001
0001
0000
0001
0002
0000
0000
0002
0000
0000
0002
0001
0001
0001
0001
0001
0000
0001
0000
0000
0001
0000
0001
0001
0000
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
0001
FFFF
0001
0001
FFFF
0002
0000
0000
0002
FFFF
0001
0001
FFFF
0001
0000
FFFF
0001
0000
0000
FFFF
0001
0001
FFFF
0000
0001
0000
0000
0001
0001
FFFF
0001
0000
FFFF
0001
0000
0000
0001
FFFF
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0001
FFFF
0000
0000
0000
0000
FFFF
0001
0000
0000
0001
FFFF
0001
0001
FFFF
0001
0000
FFFF
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFE
0001
FFFF
FFFE
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0001
0001
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0001
FFFF
0000
0001
0000
0002
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0001
0001
0000
0001
0001
0000
0001
0001
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0001
0000
0001
0001
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0001
0000
0001
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0001
0000
0000
0001
FFFF
0001
0001
FFFF
0002
0001
FFFF
0001
0000
0001
0000
FFFF
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0001
FFFF
0001
0001
FFFF
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0001
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0001
0000
0001
0002
0000
0001
0001
FFFF
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0001
0001
0000
0001
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0001
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
0000
FFFE
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
0002
0000
FFFF
0001
FFFF
0000
0001
0000
0000
0001
0001
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0001
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0001
0000
0000
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFE
0000
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
FFFF
0000
0001
0000
0000
0000
0000
FFFF
0000
0002
0000
0000
0001
FFFF
0000
0000
FFFF
0001
0000
0000
FFFF
0000
0001
FFFF
FFFF
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0001
0001
0000
0000
0001
0001
0000
0001
0001
FFFF
0001
0001
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0001
FFFF
0001
0000
FFFF
0002
FFFF
FFFF
0001
FFFF
0000
FFFF
0000
0000
FFFE
0001
0000
FFFF
0001
FFFF
0001
0000
FFFF
0001
0000
FFFF
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0001
0000
0000
0001
FFFF
0001
0000
FFFF
0001
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFE
0000
FFFF
FFFF
0000
FFFF
0001
0001
0000
0001
0000
0000
0001
0000
0001
0000
0000
0001
0001
0001
0000
0001
0002
0001
0000
0001
0001
0000
0001
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
0000
0000
FFFE
0001
0000
FFFE
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0001
0000
0000
0001
0000
0001
0001
FFFF
0000
0001
FFFF
0000
0001
FFFF
0001
FFFF
FFFF
0001
FFFF
0000
0001
FFFE
0001
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
FFFF
0000
0001
FFFF
0001
0000
FFFF
0002
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0001
0000
0000
0001
FFFF
0001
0001
FFFF
0001
0001
FFFF
0001
0000
0000
0001
0000
0001
0000
0001
0001
0000
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0001
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
FFFF
FFFF
0001
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0002
FFFF
FFFF
0001
FFFF
0000
0000
FFFE
0000
0000
FFFF
0001
FFFF
FFFF
0000
FFFF
0000
0001
FFFF
FFFF
0001
0000
0000
0000
0000
0001
0000
0001
0001
FFFF
0001
0001
FFFF
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
FFFF
0001
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0001
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0001
0000
FFFF
0001
FFFF
FFFF
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0001
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
0001
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0001
0001
0000
0001
0000
0001
0001
0000
0002
0000
0000
0002
FFFF
0001
0001
FFFF
0001
0001
0000
0001
0001
0001
0001
0001
0001
0000
0001
0001
0000
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0001
0000
0000
0001
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0000
0000
0001
0000
0000
0001
0001
0000
0001
0002
0000
0000
0001
0000
0000
0000
FFFF
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0001
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
0000
FFFF
0000
0000
0000
FFFF
0000
FFFF
0000
0001
0000
0000
0001
0001
0001
0000
0001
0001
0000
0001
0000
0000
0001
0000
0000
0001
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
FFFF
0001
0001
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
FFFF
0001
0001
0000
0001
0001
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0001
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0002
0000
FFFF
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0001
FFFF
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0001
FFFF
0000
0001
FFFE
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
0001
FFFF
FFFF
0001
0000
0000
0000
0001
0001
FFFF
0000
0001
0000
0000
0001
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0001
0001
0001
0000
0001
0000
0001
0000
FFFF
0002
0000
0001
0002
0000
0001
0002
0001
0001
0001
0001
0001
0001
0002
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0001
0001
0000
0001
0001
0000
0001
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0000
FFFF
0001
0000
0000
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
0000
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0001
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
0000
0001
FFFF
0002
0000
FFFF
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0000
0000
0000
0001
0001
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
FFFF
0000
0001
FFFF
0002
0000
FFFF
0001
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0001
0000
FFFF
0001
0000
0000
0001
FFFF
FFFF
0001
FFFF
0000
FFFF
FFFF
0001
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
0001
FFFF
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0000
0001
0000
FFFF
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0000
0001
0001
FFFF
0001
0001
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0002
0001
0001
0001
0001
0002
0001
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0000
0000
0001
0000
0001
0001
FFFF
0001
0001
0000
0000
0001
0001
FFFF
0000
0001
FFFF
0001
0000
FFFF
0001
FFFF
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
FFFF
0000
0001
FFFF
0000
0000
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
0001
0000
0000
0001
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0001
0000
0000
0001
0000
0001
0000
FFFF
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0001
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
0001
FFFF
0000
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0001
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0001
0001
0001
0000
0001
0001
FFFF
0001
0001
FFFF
0001
0000
0000
0001
0000
0001
0001
0000
0001
0001
0000
0000
0002
0001
0000
0002
0001
0000
0002
0000
0000
0002
FFFF
0000
0001
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0001
0000
0001
0000
0000
0001
0000
0000
0000
FFFF
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0000
0001
0000
0000
0001
FFFF
0000
0001
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
FFFF
0001
0000
FFFF
0001
0000
FFFF
0001
FFFF
FFFF
0001
FFFF
FFFF
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
FFFF
FFFF
0001
FFFF
FFFF
0000
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
FFFF
FFFE
0000
FFFF
FFFE
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
0000
0000
FFFE
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0000
FFFF
0001
0000
0000
0001
0000
0001
0002
0001
0000
0001
0002
0001
0000
0001
0001
0000
0000
0002
0000
0001
0002
0000
0000
0001
0000
0000
0000
FFFF
0001
0001
FFFF
0001
0001
0000
0001
0001
0001
0000
0001
0001
0000
0001
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0001
0001
0000
0001
0000
0001
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
0000
0000
FFFF
FFFF
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0001
0000
FFFF
0001
0001
FFFF
0001
0000
0000
0001
FFFF
FFFF
0001
FFFF
FFFF
0001
0000
FFFF
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0001
0001
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
FFFF
0000
0001
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFF
0000
0001
0000
0000
0000
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
FFFE
0000
0000
FFFE
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFE
0000
0000
FFFE
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0001
0001
0002
0001
0000
0002
0001
0000
0001
0001
0002
0000
0001
0002
0001
0001
0000
0001
0000
0000
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0000
0001
0001
0000
0001
0000
0000
0001
0000
0000
0001
0000
0000
0001
0001
0001
0000
0000
0002
FFFF
0001
0001
FFFF
0000
0000
0000
0000
0000
0001
0000
0001
0001
FFFF
0002
0000
FFFF
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
FFFF
FFFF
0000
FFFF
0000
FFFF
0000
0000
FFFE
0001
0000
FFFF
0001
FFFF
FFFF
0000
FFFF
0000
0000
0000
0001
FFFF
0000
0001
FFFF
0001
0000
0000
0001
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
FFFE
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFE
FFFF
0000
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0001
0001
FFFF
0001
0001
FFFF
0001
0000
0000
0001
0000
FFFF
0001
0000
FFFF
0001
0000
0000
0001
FFFF
0001
0001
FFFF
0001
0000
0000
0002
0000
0001
0001
0000
0002
0000
0000
0001
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0001
0000
0000
0001
0000
FFFF
0000
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
FFFF
0002
0001
0000
0001
0000
0000
0001
0000
0001
0000
FFFF
0000
FFFF
FFFF
0000
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
FFFF
0000
0001
0001
0001
0000
0001
0001
0000
0001
0000
0000
0001
FFFF
0000
0000
FFFF
0001
0000
FFFF
0000
0000
FFFF
0000
0001
FFFF
FFFF
0001
0000
0000
0001
0000
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
