2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h1 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h2 2'h2 2'h2 2'h2 2'h1 2'h2 2'h2 2'h2 2'h2 2'h1 2'h0 2'h0 2'h0
2'h0 2'h0 2'h1 2'h3 2'h3 2'h2 2'h2 2'h1 2'h3 2'h3 2'h2 2'h2 2'h1 2'h0 2'h0 2'h0
2'h0 2'h1 2'h1 2'h3 2'h3 2'h2 2'h2 2'h1 2'h3 2'h3 2'h2 2'h2 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h2 2'h2 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h1 2'h0 2'h0
2'h0 2'h1 2'h1 2'h0 2'h1 2'h1 2'h1 2'h0 2'h0 2'h1 2'h1 2'h1 2'h0 2'h1 2'h1 2'h0
2'h0 2'h1 2'h0 2'h0 2'h0 2'h1 2'h1 2'h0 2'h0 2'h1 2'h1 2'h0 2'h0 2'h0 2'h1 2'h0
2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0 2'h0

0000000000000000
0000001111000000
0000111111110000
0001331113311000
0012332123321100
0012222122221100
0012222122221100
0111221112211110
0111111111111110
0111111111111110
0111111111111110
0111111111111110
0111111111111110
0110111001110110
0100011001100010
0000000000000000
