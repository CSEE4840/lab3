// characters.vh
// 8x16 bitmap font for A-Z and 0-9

localparam logic [7:0] char_bitmaps [0:35][0:15] = '{
    // A (index 0)
    '{8'h18, 8'h3C, 8'h66, 8'hC3, 8'hC3, 8'hFF, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // B
    '{8'hFE, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h66, 8'h66, 8'h66, 8'h66, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // C
    '{8'h3C, 8'h66, 8'hC2, 8'hC0, 8'hC0, 8'hC0, 8'hC0, 8'hC2, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // D
    '{8'hFC, 8'h66, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h66, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // E
    '{8'hFF, 8'h63, 8'h68, 8'h68, 8'h78, 8'h68, 8'h68, 8'h60, 8'h63, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // F
    '{8'hFF, 8'h63, 8'h68, 8'h68, 8'h78, 8'h68, 8'h68, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // G
    '{8'h3C, 8'h66, 8'hC2, 8'hC0, 8'hC0, 8'hCF, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // H
    '{8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hFF, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // I
    '{8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // J
    '{8'h1F, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'hCC, 8'hCC, 8'h78, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // K
    '{8'hE7, 8'h66, 8'h6C, 8'h78, 8'h70, 8'h78, 8'h6C, 8'h66, 8'h66, 8'hE7, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // L
    '{8'hF0, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h63, 8'h63, 8'h63, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // M
    '{8'hC3, 8'hE7, 8'hFF, 8'hDB, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // N
    '{8'hC3, 8'hE3, 8'hF3, 8'hDB, 8'hCF, 8'hC7, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // O
    '{8'h3C, 8'h66, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // P
    '{8'hFE, 8'h66, 8'h66, 8'h66, 8'h7E, 8'h60, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // Q
    '{8'h3C, 8'h66, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hCB, 8'hC7, 8'h66, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // R
    '{8'hFE, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h78, 8'h6C, 8'h66, 8'h66, 8'hE7, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // S
    '{8'h3E, 8'h66, 8'hC0, 8'hC0, 8'h7C, 8'h06, 8'h03, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // T
    '{8'hFF, 8'hDB, 8'h99, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // U
    '{8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // V
    '{8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // W
    '{8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hDB, 8'hFF, 8'hE7, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // X
    '{8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h3C, 8'h66, 8'hC3, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // Y
    '{8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // Z
    '{8'hFF, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC0, 8'hC0, 8'hC3, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},

    // 0 (index 26)
    '{8'h3C, 8'h66, 8'hC3, 8'hC7, 8'hCF, 8'hDB, 8'hE3, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 1
    '{8'h18, 8'h38, 8'h78, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 2
    '{8'h3C, 8'h66, 8'hC3, 8'h03, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 3
    '{8'h3C, 8'h66, 8'hC3, 8'h03, 8'h1E, 8'h03, 8'h03, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 4
    '{8'h06, 8'h0E, 8'h1E, 8'h36, 8'h66, 8'hFF, 8'h06, 8'h06, 8'h06, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 5
    '{8'hFF, 8'hC0, 8'hC0, 8'hFC, 8'h06, 8'h03, 8'h03, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 6
    '{8'h3C, 8'h66, 8'hC0, 8'hC0, 8'hFC, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 7
    '{8'hFF, 8'h03, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h60, 8'h60, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 8
    '{8'h3C, 8'h66, 8'hC3, 8'h66, 8'h3C, 8'h66, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
    // 9
    '{8'h3C, 8'h66, 8'hC3, 8'hC3, 8'h67, 8'h3F, 8'h03, 8'h03, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}
};
