00000000
00003C00
00FFFF00
03FFFFC0
114719DC
1CBAAE1C
1DCECE1C
73CECE7E
74719DFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
6E1C3B1A
43198642
00000000
