00000000
00003C00
00FFFF00
04F33CC0
13B29CE4
1CAAAB9C
1CAAAB9C
74719DFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
7FFFFFFE
6E1C3B1A
43198642
00000000
